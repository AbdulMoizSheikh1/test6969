magic
tech gf180mcuD
magscale 1 5
timestamp 1701944771
<< metal2 >>
rect 5516 297780 5628 298500
rect 16548 297780 16660 298500
rect 27580 297780 27692 298500
rect 38612 297780 38724 298500
rect 49644 297780 49756 298500
rect 60676 297780 60788 298500
rect 71708 297780 71820 298500
rect 82740 297780 82852 298500
rect 93772 297780 93884 298500
rect 104804 297780 104916 298500
rect 115836 297780 115948 298500
rect 126868 297780 126980 298500
rect 137900 297780 138012 298500
rect 148932 297780 149044 298500
rect 159964 297780 160076 298500
rect 170996 297780 171108 298500
rect 182028 297780 182140 298500
rect 193060 297780 193172 298500
rect 204092 297780 204204 298500
rect 215124 297780 215236 298500
rect 226156 297780 226268 298500
rect 237188 297780 237300 298500
rect 248220 297780 248332 298500
rect 259252 297780 259364 298500
rect 270284 297780 270396 298500
rect 281316 297780 281428 298500
rect 292348 297780 292460 298500
rect 98686 238042 98714 238047
rect 98686 131306 98714 238014
rect 281414 156338 281442 156343
rect 281414 155554 281442 156310
rect 281414 155521 281442 155526
rect 98686 131273 98714 131278
rect 281470 126882 281498 126887
rect 281470 122514 281498 126854
rect 281470 122481 281498 122486
rect 282142 119322 282170 119327
rect 282142 102690 282170 119294
rect 282142 102657 282170 102662
rect 282198 104930 282226 104935
rect 104566 98938 104594 98943
rect 96166 98826 96194 98831
rect 58366 98770 58394 98775
rect 5670 98714 5698 98719
rect 5670 240 5698 98686
rect 11382 97874 11410 97879
rect 6622 27314 6650 27319
rect 6622 240 6650 27286
rect 7574 9674 7602 9679
rect 7574 240 7602 9646
rect 8638 3794 8666 3799
rect 8638 240 8666 3766
rect 10542 2170 10570 2175
rect 9590 2114 9618 2119
rect 9590 240 9618 2086
rect 10542 240 10570 2142
rect 5670 196 5796 240
rect 6622 196 6748 240
rect 7574 196 7700 240
rect 5684 -480 5796 196
rect 6636 -480 6748 196
rect 7588 -480 7700 196
rect 8540 196 8666 240
rect 9492 196 9618 240
rect 10444 196 10570 240
rect 11382 240 11410 97846
rect 15190 97034 15218 97039
rect 14294 61754 14322 61759
rect 13398 4634 13426 4639
rect 12446 3850 12474 3855
rect 12446 240 12474 3822
rect 13398 240 13426 4606
rect 14294 240 14322 61726
rect 15190 240 15218 97006
rect 43750 96194 43778 96199
rect 24710 86954 24738 86959
rect 17094 84434 17122 84439
rect 16254 4690 16282 4695
rect 16254 240 16282 4662
rect 11382 196 11508 240
rect 8540 -480 8652 196
rect 9492 -480 9604 196
rect 10444 -480 10556 196
rect 11396 -480 11508 196
rect 12348 196 12474 240
rect 13300 196 13426 240
rect 12348 -480 12460 196
rect 13300 -480 13412 196
rect 14252 -480 14364 240
rect 15190 196 15316 240
rect 15204 -480 15316 196
rect 16156 196 16282 240
rect 17094 240 17122 84406
rect 21406 81074 21434 81079
rect 18998 54194 19026 54199
rect 18158 2226 18186 2231
rect 18158 240 18186 2198
rect 17094 196 17220 240
rect 16156 -480 16268 196
rect 17108 -480 17220 196
rect 18060 196 18186 240
rect 18998 240 19026 54166
rect 20902 14714 20930 14719
rect 20062 2058 20090 2063
rect 20062 240 20090 2030
rect 18998 196 19124 240
rect 18060 -480 18172 196
rect 19012 -480 19124 196
rect 19964 196 20090 240
rect 20902 240 20930 14686
rect 21406 2058 21434 81046
rect 22806 80234 22834 80239
rect 21406 2025 21434 2030
rect 21966 2282 21994 2287
rect 21966 240 21994 2254
rect 20902 196 21028 240
rect 19964 -480 20076 196
rect 20916 -480 21028 196
rect 21868 196 21994 240
rect 22806 240 22834 80206
rect 23758 52514 23786 52519
rect 23758 240 23786 52486
rect 24710 240 24738 86926
rect 26614 79394 26642 79399
rect 25774 2338 25802 2343
rect 25774 240 25802 2310
rect 22806 196 22932 240
rect 23758 196 23884 240
rect 24710 196 24836 240
rect 21868 -480 21980 196
rect 22820 -480 22932 196
rect 23772 -480 23884 196
rect 24724 -480 24836 196
rect 25676 196 25802 240
rect 26614 240 26642 79366
rect 29470 78554 29498 78559
rect 28574 28154 28602 28159
rect 27566 26474 27594 26479
rect 27566 240 27594 26446
rect 28574 240 28602 28126
rect 29470 240 29498 78526
rect 32326 77714 32354 77719
rect 31374 42434 31402 42439
rect 30422 33194 30450 33199
rect 30422 240 30450 33166
rect 31374 240 31402 42406
rect 32326 240 32354 77686
rect 35182 76034 35210 76039
rect 34230 15554 34258 15559
rect 33390 5474 33418 5479
rect 33390 240 33418 5446
rect 26614 196 26740 240
rect 27566 196 27692 240
rect 25676 -480 25788 196
rect 26628 -480 26740 196
rect 27580 -480 27692 196
rect 28532 -480 28644 240
rect 29470 196 29596 240
rect 30422 196 30548 240
rect 31374 196 31500 240
rect 32326 196 32452 240
rect 29484 -480 29596 196
rect 30436 -480 30548 196
rect 31388 -480 31500 196
rect 32340 -480 32452 196
rect 33292 196 33418 240
rect 34230 240 34258 15526
rect 35182 240 35210 76006
rect 38038 75194 38066 75199
rect 37086 48314 37114 48319
rect 36134 6314 36162 6319
rect 36134 240 36162 6286
rect 37086 240 37114 48286
rect 38038 240 38066 75166
rect 39942 66794 39970 66799
rect 38990 6370 39018 6375
rect 38990 240 39018 6342
rect 39942 240 39970 66766
rect 42854 64274 42882 64279
rect 41846 7154 41874 7159
rect 41006 3906 41034 3911
rect 41006 240 41034 3878
rect 34230 196 34356 240
rect 35182 196 35308 240
rect 36134 196 36260 240
rect 37086 196 37212 240
rect 38038 196 38164 240
rect 38990 196 39116 240
rect 39942 196 40068 240
rect 33292 -480 33404 196
rect 34244 -480 34356 196
rect 35196 -480 35308 196
rect 36148 -480 36260 196
rect 37100 -480 37212 196
rect 38052 -480 38164 196
rect 39004 -480 39116 196
rect 39956 -480 40068 196
rect 40908 196 41034 240
rect 41846 240 41874 7126
rect 42854 240 42882 64246
rect 43750 240 43778 96166
rect 46606 93674 46634 93679
rect 44702 34034 44730 34039
rect 44702 240 44730 34006
rect 45654 7210 45682 7215
rect 45654 240 45682 7182
rect 46606 240 46634 93646
rect 52318 92834 52346 92839
rect 51366 58394 51394 58399
rect 47558 55034 47586 55039
rect 47558 240 47586 55006
rect 48510 43274 48538 43279
rect 48510 240 48538 43246
rect 50414 13034 50442 13039
rect 49518 3010 49546 3015
rect 49518 240 49546 2982
rect 50414 240 50442 13006
rect 51366 240 51394 58366
rect 52318 240 52346 92806
rect 55174 91154 55202 91159
rect 53270 34874 53298 34879
rect 53270 240 53298 34846
rect 54222 7994 54250 7999
rect 54222 240 54250 7966
rect 55174 240 55202 91126
rect 56126 56714 56154 56719
rect 56126 240 56154 56686
rect 57134 8050 57162 8055
rect 57134 240 57162 8022
rect 58366 3010 58394 98742
rect 86590 97930 86618 97935
rect 68502 97090 68530 97095
rect 66598 90314 66626 90319
rect 64694 72674 64722 72679
rect 62790 70154 62818 70159
rect 61838 44954 61866 44959
rect 58366 2977 58394 2982
rect 58982 30674 59010 30679
rect 58142 2954 58170 2959
rect 58142 240 58170 2926
rect 41846 196 41972 240
rect 40908 -480 41020 196
rect 41860 -480 41972 196
rect 42812 -480 42924 240
rect 43750 196 43876 240
rect 44702 196 44828 240
rect 45654 196 45780 240
rect 46606 196 46732 240
rect 47558 196 47684 240
rect 48510 196 48636 240
rect 43764 -480 43876 196
rect 44716 -480 44828 196
rect 45668 -480 45780 196
rect 46620 -480 46732 196
rect 47572 -480 47684 196
rect 48524 -480 48636 196
rect 49476 -480 49588 240
rect 50414 196 50540 240
rect 51366 196 51492 240
rect 52318 196 52444 240
rect 53270 196 53396 240
rect 54222 196 54348 240
rect 55174 196 55300 240
rect 56126 196 56252 240
rect 50428 -480 50540 196
rect 51380 -480 51492 196
rect 52332 -480 52444 196
rect 53284 -480 53396 196
rect 54236 -480 54348 196
rect 55188 -480 55300 196
rect 56140 -480 56252 196
rect 57092 -480 57204 240
rect 58044 196 58170 240
rect 58982 240 59010 30646
rect 59934 8106 59962 8111
rect 59934 240 59962 8078
rect 60998 3010 61026 3015
rect 60998 240 61026 2982
rect 58982 196 59108 240
rect 59934 196 60060 240
rect 58044 -480 58156 196
rect 58996 -480 59108 196
rect 59948 -480 60060 196
rect 60900 196 61026 240
rect 61838 240 61866 44926
rect 62790 240 62818 70126
rect 63798 3066 63826 3071
rect 63798 240 63826 3038
rect 64694 240 64722 72646
rect 65646 12194 65674 12199
rect 65646 240 65674 12166
rect 66598 240 66626 90286
rect 67550 57554 67578 57559
rect 67550 240 67578 57526
rect 68502 240 68530 97062
rect 69454 89474 69482 89479
rect 69454 240 69482 89446
rect 72310 87794 72338 87799
rect 71414 8834 71442 8839
rect 70406 6426 70434 6431
rect 70406 240 70434 6398
rect 71414 240 71442 8806
rect 72310 240 72338 87766
rect 75166 87010 75194 87015
rect 73262 71834 73290 71839
rect 73262 240 73290 71806
rect 74214 8890 74242 8895
rect 74214 240 74242 8862
rect 75166 240 75194 86982
rect 78022 85274 78050 85279
rect 76118 70994 76146 70999
rect 76118 240 76146 70966
rect 77070 37394 77098 37399
rect 77070 240 77098 37366
rect 78022 240 78050 85246
rect 83734 84490 83762 84495
rect 82782 53354 82810 53359
rect 81830 18914 81858 18919
rect 80878 12250 80906 12255
rect 78974 9730 79002 9735
rect 78974 240 79002 9702
rect 79926 8946 79954 8951
rect 79926 240 79954 8918
rect 80878 240 80906 12222
rect 81830 240 81858 18886
rect 82782 240 82810 53326
rect 83734 240 83762 84462
rect 85694 44114 85722 44119
rect 84686 7266 84714 7271
rect 84686 240 84714 7238
rect 85694 240 85722 44086
rect 86590 240 86618 97902
rect 91350 92890 91378 92895
rect 89446 88634 89474 88639
rect 87542 65954 87570 65959
rect 87542 240 87570 65926
rect 88494 60074 88522 60079
rect 88494 240 88522 60046
rect 89446 240 89474 88606
rect 90398 36554 90426 36559
rect 90398 240 90426 36526
rect 91350 240 91378 92862
rect 94206 91210 94234 91215
rect 92302 81130 92330 81135
rect 92302 240 92330 81102
rect 93254 51674 93282 51679
rect 93254 240 93282 51646
rect 94206 240 94234 91182
rect 96110 22274 96138 22279
rect 95270 2562 95298 2567
rect 95270 240 95298 2534
rect 61838 196 61964 240
rect 62790 196 62916 240
rect 60900 -480 61012 196
rect 61852 -480 61964 196
rect 62804 -480 62916 196
rect 63756 -480 63868 240
rect 64694 196 64820 240
rect 65646 196 65772 240
rect 66598 196 66724 240
rect 67550 196 67676 240
rect 68502 196 68628 240
rect 69454 196 69580 240
rect 70406 196 70532 240
rect 64708 -480 64820 196
rect 65660 -480 65772 196
rect 66612 -480 66724 196
rect 67564 -480 67676 196
rect 68516 -480 68628 196
rect 69468 -480 69580 196
rect 70420 -480 70532 196
rect 71372 -480 71484 240
rect 72310 196 72436 240
rect 73262 196 73388 240
rect 74214 196 74340 240
rect 75166 196 75292 240
rect 76118 196 76244 240
rect 77070 196 77196 240
rect 78022 196 78148 240
rect 78974 196 79100 240
rect 79926 196 80052 240
rect 80878 196 81004 240
rect 81830 196 81956 240
rect 82782 196 82908 240
rect 83734 196 83860 240
rect 84686 196 84812 240
rect 72324 -480 72436 196
rect 73276 -480 73388 196
rect 74228 -480 74340 196
rect 75180 -480 75292 196
rect 76132 -480 76244 196
rect 77084 -480 77196 196
rect 78036 -480 78148 196
rect 78988 -480 79100 196
rect 79940 -480 80052 196
rect 80892 -480 81004 196
rect 81844 -480 81956 196
rect 82796 -480 82908 196
rect 83748 -480 83860 196
rect 84700 -480 84812 196
rect 85652 -480 85764 240
rect 86590 196 86716 240
rect 87542 196 87668 240
rect 88494 196 88620 240
rect 89446 196 89572 240
rect 90398 196 90524 240
rect 91350 196 91476 240
rect 92302 196 92428 240
rect 93254 196 93380 240
rect 94206 196 94332 240
rect 86604 -480 86716 196
rect 87556 -480 87668 196
rect 88508 -480 88620 196
rect 89460 -480 89572 196
rect 90412 -480 90524 196
rect 91364 -480 91476 196
rect 92316 -480 92428 196
rect 93268 -480 93380 196
rect 94220 -480 94332 196
rect 95172 196 95298 240
rect 96110 240 96138 22246
rect 96166 2562 96194 98798
rect 96166 2529 96194 2534
rect 98014 96250 98042 96255
rect 97174 1274 97202 1279
rect 97174 240 97202 1246
rect 96110 196 96236 240
rect 95172 -480 95284 196
rect 96124 -480 96236 196
rect 97076 196 97202 240
rect 98014 240 98042 96222
rect 103726 93730 103754 93735
rect 100870 81914 100898 81919
rect 99974 39074 100002 39079
rect 98966 18074 98994 18079
rect 98966 240 98994 18046
rect 99974 240 100002 39046
rect 100870 240 100898 81886
rect 101822 69314 101850 69319
rect 101822 240 101850 69286
rect 102774 39914 102802 39919
rect 102774 240 102802 39886
rect 103726 240 103754 93702
rect 104566 12250 104594 98910
rect 105798 98882 105826 98887
rect 104566 12217 104594 12222
rect 104678 35714 104706 35719
rect 104678 240 104706 35686
rect 105630 21434 105658 21439
rect 105630 240 105658 21406
rect 105798 2562 105826 98854
rect 105966 98714 105994 100044
rect 105966 98681 105994 98686
rect 106526 27314 106554 100044
rect 106526 27281 106554 27286
rect 107086 9674 107114 100044
rect 107086 9641 107114 9646
rect 107534 9674 107562 9679
rect 105798 2529 105826 2534
rect 106582 2562 106610 2567
rect 106582 240 106610 2534
rect 107534 240 107562 9646
rect 107646 3794 107674 100044
rect 107646 3761 107674 3766
rect 108206 2114 108234 100044
rect 108206 2081 108234 2086
rect 108486 29834 108514 29839
rect 108486 240 108514 29806
rect 108766 2170 108794 100044
rect 109326 97874 109354 100044
rect 109326 97841 109354 97846
rect 108766 2137 108794 2142
rect 109438 13090 109466 13095
rect 109438 240 109466 13062
rect 109886 3850 109914 100044
rect 110446 4634 110474 100044
rect 111006 61754 111034 100044
rect 111566 97034 111594 100044
rect 111566 97001 111594 97006
rect 111006 61721 111034 61726
rect 111342 24794 111370 24799
rect 110446 4601 110474 4606
rect 110502 4746 110530 4751
rect 109886 3817 109914 3822
rect 110502 240 110530 4718
rect 98014 196 98140 240
rect 98966 196 99092 240
rect 97076 -480 97188 196
rect 98028 -480 98140 196
rect 98980 -480 99092 196
rect 99932 -480 100044 240
rect 100870 196 100996 240
rect 101822 196 101948 240
rect 102774 196 102900 240
rect 103726 196 103852 240
rect 104678 196 104804 240
rect 105630 196 105756 240
rect 106582 196 106708 240
rect 107534 196 107660 240
rect 108486 196 108612 240
rect 109438 196 109564 240
rect 100884 -480 100996 196
rect 101836 -480 101948 196
rect 102788 -480 102900 196
rect 103740 -480 103852 196
rect 104692 -480 104804 196
rect 105644 -480 105756 196
rect 106596 -480 106708 196
rect 107548 -480 107660 196
rect 108500 -480 108612 196
rect 109452 -480 109564 196
rect 110404 196 110530 240
rect 111342 240 111370 24766
rect 112126 4690 112154 100044
rect 112686 84434 112714 100044
rect 112686 84401 112714 84406
rect 112126 4657 112154 4662
rect 112406 3794 112434 3799
rect 112406 240 112434 3766
rect 113246 2226 113274 100044
rect 113806 54194 113834 100044
rect 114366 81074 114394 100044
rect 114366 81041 114394 81046
rect 113806 54161 113834 54166
rect 114254 23954 114282 23959
rect 113246 2193 113274 2198
rect 113302 16394 113330 16399
rect 113302 240 113330 16366
rect 114254 240 114282 23926
rect 114926 14714 114954 100044
rect 114926 14681 114954 14686
rect 115150 14714 115178 14719
rect 115150 240 115178 14686
rect 115486 2282 115514 100044
rect 116046 80234 116074 100044
rect 116046 80201 116074 80206
rect 116606 52514 116634 100044
rect 116606 52481 116634 52486
rect 117054 97034 117082 97039
rect 115486 2249 115514 2254
rect 116102 25634 116130 25639
rect 116102 240 116130 25606
rect 117054 240 117082 97006
rect 117166 86954 117194 100044
rect 117166 86921 117194 86926
rect 117726 2338 117754 100044
rect 118286 79394 118314 100044
rect 118286 79361 118314 79366
rect 118846 26474 118874 100044
rect 119406 28154 119434 100044
rect 119966 78554 119994 100044
rect 119966 78521 119994 78526
rect 120526 33194 120554 100044
rect 121086 42434 121114 100044
rect 121646 77714 121674 100044
rect 121646 77681 121674 77686
rect 121086 42401 121114 42406
rect 120526 33161 120554 33166
rect 119406 28121 119434 28126
rect 121814 27314 121842 27319
rect 118846 26441 118874 26446
rect 118958 26474 118986 26479
rect 117726 2305 117754 2310
rect 118006 12250 118034 12255
rect 118006 240 118034 12222
rect 118958 240 118986 26446
rect 119910 17290 119938 17295
rect 119910 240 119938 17262
rect 120862 15610 120890 15615
rect 120862 240 120890 15582
rect 121814 240 121842 27286
rect 122206 5474 122234 100044
rect 122766 15554 122794 100044
rect 123326 76034 123354 100044
rect 123326 76001 123354 76006
rect 122766 15521 122794 15526
rect 123718 17234 123746 17239
rect 122206 5441 122234 5446
rect 122878 3850 122906 3855
rect 122878 240 122906 3822
rect 111342 196 111468 240
rect 110404 -480 110516 196
rect 111356 -480 111468 196
rect 112308 196 112434 240
rect 112308 -480 112420 196
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115150 196 115276 240
rect 116102 196 116228 240
rect 117054 196 117180 240
rect 118006 196 118132 240
rect 118958 196 119084 240
rect 119910 196 120036 240
rect 120862 196 120988 240
rect 121814 196 121940 240
rect 115164 -480 115276 196
rect 116116 -480 116228 196
rect 117068 -480 117180 196
rect 118020 -480 118132 196
rect 118972 -480 119084 196
rect 119924 -480 120036 196
rect 120876 -480 120988 196
rect 121828 -480 121940 196
rect 122780 196 122906 240
rect 123718 240 123746 17206
rect 123886 6314 123914 100044
rect 124278 98322 124306 98327
rect 124278 96194 124306 98294
rect 124278 96161 124306 96166
rect 124446 48314 124474 100044
rect 125006 75194 125034 100044
rect 125006 75161 125034 75166
rect 124446 48281 124474 48286
rect 123886 6281 123914 6286
rect 124670 10514 124698 10519
rect 124670 240 124698 10486
rect 125566 6370 125594 100044
rect 126126 66794 126154 100044
rect 126126 66761 126154 66766
rect 125566 6337 125594 6342
rect 126574 18130 126602 18135
rect 125734 4634 125762 4639
rect 125734 240 125762 4606
rect 123718 196 123844 240
rect 124670 196 124796 240
rect 122780 -480 122892 196
rect 123732 -480 123844 196
rect 124684 -480 124796 196
rect 125636 196 125762 240
rect 126574 240 126602 18102
rect 126686 3906 126714 100044
rect 127246 7154 127274 100044
rect 127806 64274 127834 100044
rect 128366 98322 128394 100044
rect 128366 98289 128394 98294
rect 127806 64241 127834 64246
rect 127246 7121 127274 7126
rect 128534 34090 128562 34095
rect 126686 3873 126714 3878
rect 127526 6314 127554 6319
rect 127526 240 127554 6286
rect 128534 240 128562 34062
rect 128926 34034 128954 100044
rect 128926 34001 128954 34006
rect 129430 18970 129458 18975
rect 129430 240 129458 18942
rect 129486 7210 129514 100044
rect 130046 93674 130074 100044
rect 130046 93641 130074 93646
rect 130606 55034 130634 100044
rect 130606 55001 130634 55006
rect 131166 43274 131194 100044
rect 131726 98770 131754 100044
rect 131726 98737 131754 98742
rect 131166 43241 131194 43246
rect 129486 7177 129514 7182
rect 130382 28154 130410 28159
rect 130382 240 130410 28126
rect 131334 16450 131362 16455
rect 131334 240 131362 16422
rect 132286 13034 132314 100044
rect 132846 58394 132874 100044
rect 133406 92834 133434 100044
rect 133406 92801 133434 92806
rect 132846 58361 132874 58366
rect 133966 34874 133994 100044
rect 133966 34841 133994 34846
rect 134190 33194 134218 33199
rect 132286 13001 132314 13006
rect 132342 21490 132370 21495
rect 132342 240 132370 21462
rect 133238 15554 133266 15559
rect 133238 240 133266 15526
rect 134190 240 134218 33166
rect 134526 7994 134554 100044
rect 135086 91154 135114 100044
rect 135086 91121 135114 91126
rect 135646 56714 135674 100044
rect 135646 56681 135674 56686
rect 135702 98714 135730 98719
rect 135702 12194 135730 98686
rect 135702 12161 135730 12166
rect 136206 8050 136234 100044
rect 136206 8017 136234 8022
rect 134526 7961 134554 7966
rect 136094 7154 136122 7159
rect 135198 3906 135226 3911
rect 135198 240 135226 3878
rect 136094 240 136122 7126
rect 136766 2954 136794 100044
rect 136766 2921 136794 2926
rect 137046 30730 137074 30735
rect 137046 240 137074 30702
rect 137326 30674 137354 100044
rect 137382 98322 137410 98327
rect 137382 72674 137410 98294
rect 137382 72641 137410 72646
rect 137326 30641 137354 30646
rect 137886 8106 137914 100044
rect 137886 8073 137914 8078
rect 137998 7994 138026 7999
rect 137998 240 138026 7966
rect 138446 3010 138474 100044
rect 139006 44954 139034 100044
rect 139062 98994 139090 98999
rect 139062 90314 139090 98966
rect 139062 90281 139090 90286
rect 139566 70154 139594 100044
rect 139566 70121 139594 70126
rect 139006 44921 139034 44926
rect 138446 2977 138474 2982
rect 138950 22330 138978 22335
rect 138950 240 138978 22302
rect 140014 5474 140042 5479
rect 140014 240 140042 5446
rect 140126 3066 140154 100044
rect 140686 98322 140714 100044
rect 141246 98714 141274 100044
rect 141806 98994 141834 100044
rect 141806 98961 141834 98966
rect 141246 98681 141274 98686
rect 140686 98289 140714 98294
rect 142366 57554 142394 100044
rect 142814 100030 142940 100058
rect 142422 99106 142450 99111
rect 142422 89474 142450 99078
rect 142814 98294 142842 100030
rect 143486 99106 143514 100044
rect 143486 99073 143514 99078
rect 142758 98266 142842 98294
rect 142758 97090 142786 98266
rect 142758 97057 142786 97062
rect 142422 89441 142450 89446
rect 142366 57521 142394 57526
rect 143710 64274 143738 64279
rect 140126 3033 140154 3038
rect 141918 3066 141946 3071
rect 140966 2954 140994 2959
rect 140966 240 140994 2926
rect 141918 240 141946 3038
rect 142870 3010 142898 3015
rect 142870 240 142898 2982
rect 126574 196 126700 240
rect 127526 196 127652 240
rect 125636 -480 125748 196
rect 126588 -480 126700 196
rect 127540 -480 127652 196
rect 128492 -480 128604 240
rect 129430 196 129556 240
rect 130382 196 130508 240
rect 131334 196 131460 240
rect 129444 -480 129556 196
rect 130396 -480 130508 196
rect 131348 -480 131460 196
rect 132300 -480 132412 240
rect 133238 196 133364 240
rect 134190 196 134316 240
rect 133252 -480 133364 196
rect 134204 -480 134316 196
rect 135156 -480 135268 240
rect 136094 196 136220 240
rect 137046 196 137172 240
rect 137998 196 138124 240
rect 138950 196 139076 240
rect 136108 -480 136220 196
rect 137060 -480 137172 196
rect 138012 -480 138124 196
rect 138964 -480 139076 196
rect 139916 196 140042 240
rect 140868 196 140994 240
rect 141820 196 141946 240
rect 142772 196 142898 240
rect 143710 240 143738 64246
rect 144046 6426 144074 100044
rect 144606 8834 144634 100044
rect 145166 87794 145194 100044
rect 145166 87761 145194 87766
rect 145670 100030 145740 100058
rect 145670 71834 145698 100030
rect 145670 71801 145698 71806
rect 145726 98714 145754 98719
rect 145614 13034 145642 13039
rect 144606 8801 144634 8806
rect 144662 9002 144690 9007
rect 144046 6393 144074 6398
rect 144662 240 144690 8974
rect 145614 240 145642 13006
rect 145726 3010 145754 98686
rect 146286 8890 146314 100044
rect 146846 87010 146874 100044
rect 146846 86977 146874 86982
rect 147406 70994 147434 100044
rect 147406 70961 147434 70966
rect 147518 97874 147546 97879
rect 146286 8857 146314 8862
rect 145726 2977 145754 2982
rect 146566 6370 146594 6375
rect 146566 240 146594 6342
rect 147518 240 147546 97846
rect 147966 37394 147994 100044
rect 148526 85274 148554 100044
rect 148526 85241 148554 85246
rect 147966 37361 147994 37366
rect 148470 14770 148498 14775
rect 148470 240 148498 14742
rect 149086 9730 149114 100044
rect 149086 9697 149114 9702
rect 149422 9730 149450 9735
rect 149422 240 149450 9702
rect 149646 8946 149674 100044
rect 150206 98938 150234 100044
rect 150206 98905 150234 98910
rect 149646 8913 149674 8918
rect 150374 24010 150402 24015
rect 150374 240 150402 23982
rect 150766 18914 150794 100044
rect 151326 53354 151354 100044
rect 151886 84490 151914 100044
rect 151886 84457 151914 84462
rect 151326 53321 151354 53326
rect 150766 18881 150794 18886
rect 151326 18914 151354 18919
rect 151326 240 151354 18886
rect 152446 7266 152474 100044
rect 153006 44114 153034 100044
rect 153566 97930 153594 100044
rect 153566 97897 153594 97902
rect 154126 65954 154154 100044
rect 154182 99050 154210 99055
rect 154182 92890 154210 99022
rect 154182 92857 154210 92862
rect 154126 65921 154154 65926
rect 154182 66010 154210 66015
rect 153006 44081 153034 44086
rect 152446 7233 152474 7238
rect 153230 8050 153258 8055
rect 152278 7210 152306 7215
rect 152278 240 152306 7182
rect 153230 240 153258 8022
rect 154182 240 154210 65982
rect 154686 60074 154714 100044
rect 155246 88634 155274 100044
rect 155246 88601 155274 88606
rect 154686 60041 154714 60046
rect 155806 36554 155834 100044
rect 155862 99106 155890 99111
rect 155862 81130 155890 99078
rect 156366 99050 156394 100044
rect 156926 99106 156954 100044
rect 156926 99073 156954 99078
rect 156366 99017 156394 99022
rect 155862 81097 155890 81102
rect 157486 51674 157514 100044
rect 157934 100030 158060 100058
rect 157486 51641 157514 51646
rect 157542 99106 157570 99111
rect 155806 36521 155834 36526
rect 157094 25690 157122 25695
rect 156086 24850 156114 24855
rect 155134 8834 155162 8839
rect 155134 240 155162 8806
rect 156086 240 156114 24822
rect 157094 240 157122 25662
rect 157542 22274 157570 99078
rect 157934 98294 157962 100030
rect 158606 98826 158634 100044
rect 159166 99106 159194 100044
rect 159166 99073 159194 99078
rect 158606 98793 158634 98798
rect 157654 98266 157962 98294
rect 159166 98770 159194 98775
rect 157654 91210 157682 98266
rect 157654 91177 157682 91182
rect 157542 22241 157570 22246
rect 158942 6426 158970 6431
rect 158102 2562 158130 2567
rect 158102 240 158130 2534
rect 143710 196 143836 240
rect 144662 196 144788 240
rect 145614 196 145740 240
rect 146566 196 146692 240
rect 147518 196 147644 240
rect 148470 196 148596 240
rect 149422 196 149548 240
rect 150374 196 150500 240
rect 151326 196 151452 240
rect 152278 196 152404 240
rect 153230 196 153356 240
rect 154182 196 154308 240
rect 155134 196 155260 240
rect 156086 196 156212 240
rect 139916 -480 140028 196
rect 140868 -480 140980 196
rect 141820 -480 141932 196
rect 142772 -480 142884 196
rect 143724 -480 143836 196
rect 144676 -480 144788 196
rect 145628 -480 145740 196
rect 146580 -480 146692 196
rect 147532 -480 147644 196
rect 148484 -480 148596 196
rect 149436 -480 149548 196
rect 150388 -480 150500 196
rect 151340 -480 151452 196
rect 152292 -480 152404 196
rect 153244 -480 153356 196
rect 154196 -480 154308 196
rect 155148 -480 155260 196
rect 156100 -480 156212 196
rect 157052 -480 157164 240
rect 158004 196 158130 240
rect 158942 240 158970 6398
rect 159166 2562 159194 98742
rect 159166 2529 159194 2534
rect 159726 1274 159754 100044
rect 160286 96250 160314 100044
rect 160286 96217 160314 96222
rect 160846 18074 160874 100044
rect 161406 39074 161434 100044
rect 161966 81914 161994 100044
rect 161966 81881 161994 81886
rect 162526 69314 162554 100044
rect 162526 69281 162554 69286
rect 162750 69314 162778 69319
rect 161406 39041 161434 39046
rect 160846 18041 160874 18046
rect 160846 12194 160874 12199
rect 159726 1241 159754 1246
rect 159894 10570 159922 10575
rect 159894 240 159922 10542
rect 160846 240 160874 12166
rect 161798 9786 161826 9791
rect 161798 240 161826 9758
rect 162750 240 162778 69286
rect 163086 39914 163114 100044
rect 163646 93730 163674 100044
rect 163646 93697 163674 93702
rect 163086 39881 163114 39886
rect 164206 35714 164234 100044
rect 164206 35681 164234 35686
rect 164766 21434 164794 100044
rect 165326 98882 165354 100044
rect 165326 98849 165354 98854
rect 164766 21401 164794 21406
rect 165606 12306 165634 12311
rect 164766 4690 164794 4695
rect 163758 3066 163786 3071
rect 163758 240 163786 3038
rect 164766 240 164794 4662
rect 158942 196 159068 240
rect 159894 196 160020 240
rect 160846 196 160972 240
rect 161798 196 161924 240
rect 162750 196 162876 240
rect 158004 -480 158116 196
rect 158956 -480 159068 196
rect 159908 -480 160020 196
rect 160860 -480 160972 196
rect 161812 -480 161924 196
rect 162764 -480 162876 196
rect 163716 -480 163828 240
rect 164668 196 164794 240
rect 165606 240 165634 12278
rect 165886 9674 165914 100044
rect 165886 9641 165914 9646
rect 165942 98826 165970 98831
rect 165942 3906 165970 98798
rect 166446 29834 166474 100044
rect 166446 29801 166474 29806
rect 165942 3873 165970 3878
rect 166558 13146 166586 13151
rect 166558 240 166586 13118
rect 167006 13090 167034 100044
rect 167006 13057 167034 13062
rect 167566 4746 167594 100044
rect 168126 24794 168154 100044
rect 168126 24761 168154 24766
rect 168462 26530 168490 26535
rect 167566 4713 167594 4718
rect 167622 3906 167650 3911
rect 167622 240 167650 3878
rect 165606 196 165732 240
rect 166558 196 166684 240
rect 164668 -480 164780 196
rect 165620 -480 165732 196
rect 166572 -480 166684 196
rect 167524 196 167650 240
rect 168462 240 168490 26502
rect 168686 3794 168714 100044
rect 169246 16394 169274 100044
rect 169302 99050 169330 99055
rect 169302 17290 169330 99022
rect 169806 23954 169834 100044
rect 169806 23921 169834 23926
rect 169302 17257 169330 17262
rect 169246 16361 169274 16366
rect 169414 16394 169442 16399
rect 168686 3761 168714 3766
rect 169414 240 169442 16366
rect 170366 14714 170394 100044
rect 170926 25634 170954 100044
rect 171374 100030 171500 100058
rect 170926 25601 170954 25606
rect 170982 99106 171010 99111
rect 170366 14681 170394 14686
rect 170422 17290 170450 17295
rect 170422 240 170450 17262
rect 170982 12250 171010 99078
rect 171374 98294 171402 100030
rect 172046 99106 172074 100044
rect 172046 99073 172074 99078
rect 171318 98266 171402 98294
rect 171318 97034 171346 98266
rect 171318 97001 171346 97006
rect 172606 26474 172634 100044
rect 172606 26441 172634 26446
rect 172662 99106 172690 99111
rect 172662 15610 172690 99078
rect 173166 99050 173194 100044
rect 173726 99106 173754 100044
rect 173726 99073 173754 99078
rect 173166 99017 173194 99022
rect 172662 15577 172690 15582
rect 172718 27370 172746 27375
rect 170982 12217 171010 12222
rect 172270 14714 172298 14719
rect 171430 2114 171458 2119
rect 171430 240 171458 2086
rect 168462 196 168588 240
rect 169414 196 169540 240
rect 167524 -480 167636 196
rect 168476 -480 168588 196
rect 169428 -480 169540 196
rect 170380 -480 170492 240
rect 171332 196 171458 240
rect 172270 240 172298 14686
rect 172718 2114 172746 27342
rect 174286 27314 174314 100044
rect 174286 27281 174314 27286
rect 174342 98994 174370 98999
rect 174174 21434 174202 21439
rect 172718 2081 172746 2086
rect 173334 3794 173362 3799
rect 173334 240 173362 3766
rect 172270 196 172396 240
rect 171332 -480 171444 196
rect 172284 -480 172396 196
rect 173236 196 173362 240
rect 174174 240 174202 21406
rect 174342 6314 174370 98966
rect 174342 6281 174370 6286
rect 174846 3850 174874 100044
rect 175406 17234 175434 100044
rect 175406 17201 175434 17206
rect 175966 10514 175994 100044
rect 175966 10481 175994 10486
rect 176022 99106 176050 99111
rect 174846 3817 174874 3822
rect 175126 6314 175154 6319
rect 175126 240 175154 6286
rect 176022 4634 176050 99078
rect 176526 99106 176554 100044
rect 176526 99073 176554 99078
rect 177086 18130 177114 100044
rect 177646 98994 177674 100044
rect 177646 98961 177674 98966
rect 177646 98882 177674 98887
rect 177646 30730 177674 98854
rect 177646 30697 177674 30702
rect 177982 76034 178010 76039
rect 177086 18097 177114 18102
rect 176022 4601 176050 4606
rect 177030 17234 177058 17239
rect 176190 3850 176218 3855
rect 176190 240 176218 3822
rect 174174 196 174300 240
rect 175126 196 175252 240
rect 173236 -480 173348 196
rect 174188 -480 174300 196
rect 175140 -480 175252 196
rect 176092 196 176218 240
rect 177030 240 177058 17206
rect 177982 240 178010 76006
rect 178206 34090 178234 100044
rect 178206 34057 178234 34062
rect 178766 18970 178794 100044
rect 179326 28154 179354 100044
rect 179326 28121 179354 28126
rect 179382 99106 179410 99111
rect 178766 18937 178794 18942
rect 178934 18074 178962 18079
rect 178934 240 178962 18046
rect 179382 16450 179410 99078
rect 179886 99106 179914 100044
rect 179886 99073 179914 99078
rect 180446 21490 180474 100044
rect 180446 21457 180474 21462
rect 179382 16417 179410 16422
rect 180838 15610 180866 15615
rect 179998 2114 180026 2119
rect 179998 240 180026 2086
rect 177030 196 177156 240
rect 177982 196 178108 240
rect 178934 196 179060 240
rect 176092 -480 176204 196
rect 177044 -480 177156 196
rect 177996 -480 178108 196
rect 178948 -480 179060 196
rect 179900 196 180026 240
rect 180838 240 180866 15582
rect 181006 15554 181034 100044
rect 181566 33194 181594 100044
rect 182126 98826 182154 100044
rect 182126 98793 182154 98798
rect 181566 33161 181594 33166
rect 181006 15521 181034 15526
rect 181790 7266 181818 7271
rect 181790 240 181818 7238
rect 182686 7154 182714 100044
rect 183246 98882 183274 100044
rect 183246 98849 183274 98854
rect 183526 29834 183554 29839
rect 182686 7121 182714 7126
rect 182854 28154 182882 28159
rect 182854 4214 182882 28126
rect 182798 4186 182882 4214
rect 182798 2170 182826 4186
rect 182798 2137 182826 2142
rect 182854 2114 182882 2119
rect 182854 240 182882 2086
rect 183526 2114 183554 29806
rect 183526 2081 183554 2086
rect 183694 8106 183722 8111
rect 180838 196 180964 240
rect 181790 196 181916 240
rect 179900 -480 180012 196
rect 180852 -480 180964 196
rect 181804 -480 181916 196
rect 182756 196 182882 240
rect 183694 240 183722 8078
rect 183806 7994 183834 100044
rect 184366 22330 184394 100044
rect 184366 22297 184394 22302
rect 184422 98826 184450 98831
rect 184422 9002 184450 98798
rect 184422 8969 184450 8974
rect 183806 7961 183834 7966
rect 184646 8890 184674 8895
rect 184646 240 184674 8862
rect 184926 5474 184954 100044
rect 184926 5441 184954 5446
rect 185486 2954 185514 100044
rect 185486 2921 185514 2926
rect 185654 22274 185682 22279
rect 185654 240 185682 22246
rect 186046 3010 186074 100044
rect 186606 98714 186634 100044
rect 186606 98681 186634 98686
rect 186102 98322 186130 98327
rect 186102 64274 186130 98294
rect 187166 98322 187194 100044
rect 187726 98826 187754 100044
rect 187726 98793 187754 98798
rect 187166 98289 187194 98294
rect 187726 98714 187754 98719
rect 186102 64241 186130 64246
rect 186046 2977 186074 2982
rect 187502 9674 187530 9679
rect 186662 2562 186690 2567
rect 186662 240 186690 2534
rect 183694 196 183820 240
rect 184646 196 184772 240
rect 182756 -480 182868 196
rect 183708 -480 183820 196
rect 184660 -480 184772 196
rect 185612 -480 185724 240
rect 186564 196 186690 240
rect 187502 240 187530 9646
rect 187726 6370 187754 98686
rect 188286 13034 188314 100044
rect 188846 98714 188874 100044
rect 188846 98681 188874 98686
rect 189406 97874 189434 100044
rect 189406 97841 189434 97846
rect 189966 14770 189994 100044
rect 189966 14737 189994 14742
rect 190246 14770 190274 14775
rect 188286 13001 188314 13006
rect 187726 6337 187754 6342
rect 189518 3122 189546 3127
rect 188566 2114 188594 2119
rect 188566 240 188594 2086
rect 189518 240 189546 3094
rect 190246 2114 190274 14742
rect 190526 9730 190554 100044
rect 191086 24010 191114 100044
rect 191086 23977 191114 23982
rect 191142 98714 191170 98719
rect 190526 9697 190554 9702
rect 190246 2081 190274 2086
rect 190358 6370 190386 6375
rect 187502 196 187628 240
rect 186564 -480 186676 196
rect 187516 -480 187628 196
rect 188468 196 188594 240
rect 189420 196 189546 240
rect 190358 240 190386 6342
rect 191142 2562 191170 98686
rect 191646 18914 191674 100044
rect 191646 18881 191674 18886
rect 192206 7210 192234 100044
rect 192766 8050 192794 100044
rect 193326 66010 193354 100044
rect 193326 65977 193354 65982
rect 192766 8017 192794 8022
rect 192822 23954 192850 23959
rect 192206 7177 192234 7182
rect 191142 2529 191170 2534
rect 192318 2954 192346 2959
rect 191422 2506 191450 2511
rect 191422 240 191450 2478
rect 192318 240 192346 2926
rect 192822 2506 192850 23926
rect 193886 8834 193914 100044
rect 194446 24850 194474 100044
rect 194446 24817 194474 24822
rect 194502 98378 194530 98383
rect 193886 8801 193914 8806
rect 192822 2473 192850 2478
rect 193214 8050 193242 8055
rect 193214 240 193242 8022
rect 194502 3066 194530 98350
rect 195006 25690 195034 100044
rect 195006 25657 195034 25662
rect 195286 99106 195314 99111
rect 195286 10570 195314 99078
rect 195566 98770 195594 100044
rect 195566 98737 195594 98742
rect 195286 10537 195314 10542
rect 195342 24794 195370 24799
rect 194502 3033 194530 3038
rect 195230 3010 195258 3015
rect 194278 2114 194306 2119
rect 194278 240 194306 2086
rect 195230 240 195258 2982
rect 195342 2114 195370 24766
rect 195342 2081 195370 2086
rect 196070 18914 196098 18919
rect 190358 196 190484 240
rect 188468 -480 188580 196
rect 189420 -480 189532 196
rect 190372 -480 190484 196
rect 191324 196 191450 240
rect 191324 -480 191436 196
rect 192276 -480 192388 240
rect 193214 196 193340 240
rect 193228 -480 193340 196
rect 194180 196 194306 240
rect 195132 196 195258 240
rect 196070 240 196098 18886
rect 196126 6426 196154 100044
rect 196686 99106 196714 100044
rect 196686 99073 196714 99078
rect 196126 6393 196154 6398
rect 197022 25634 197050 25639
rect 197022 240 197050 25606
rect 197246 12194 197274 100044
rect 197246 12161 197274 12166
rect 197806 9786 197834 100044
rect 198366 69314 198394 100044
rect 198366 69281 198394 69286
rect 198646 99106 198674 99111
rect 198646 17290 198674 99078
rect 198926 98378 198954 100044
rect 198926 98345 198954 98350
rect 198646 17257 198674 17262
rect 197806 9753 197834 9758
rect 198926 12194 198954 12199
rect 197974 7154 198002 7159
rect 197974 240 198002 7126
rect 198926 240 198954 12166
rect 199486 4690 199514 100044
rect 199486 4657 199514 4662
rect 199542 98770 199570 98775
rect 199542 3122 199570 98742
rect 200046 12306 200074 100044
rect 200606 13146 200634 100044
rect 200606 13113 200634 13118
rect 200830 42434 200858 42439
rect 200046 12273 200074 12278
rect 199542 3089 199570 3094
rect 199934 10514 199962 10519
rect 199934 240 199962 10486
rect 200830 240 200858 42406
rect 201166 3906 201194 100044
rect 201726 26530 201754 100044
rect 201726 26497 201754 26502
rect 202286 16394 202314 100044
rect 202846 99106 202874 100044
rect 202846 99073 202874 99078
rect 203406 27370 203434 100044
rect 203406 27337 203434 27342
rect 202286 16361 202314 16366
rect 203742 16394 203770 16399
rect 201166 3873 201194 3878
rect 201782 13034 201810 13039
rect 201782 240 201810 13006
rect 203686 8834 203714 8839
rect 202846 2114 202874 2119
rect 202846 240 202874 2086
rect 196070 196 196196 240
rect 197022 196 197148 240
rect 197974 196 198100 240
rect 198926 196 199052 240
rect 194180 -480 194292 196
rect 195132 -480 195244 196
rect 196084 -480 196196 196
rect 197036 -480 197148 196
rect 197988 -480 198100 196
rect 198940 -480 199052 196
rect 199892 -480 200004 240
rect 200830 196 200956 240
rect 201782 196 201908 240
rect 200844 -480 200956 196
rect 201796 -480 201908 196
rect 202748 196 202874 240
rect 203686 240 203714 8806
rect 203742 2114 203770 16366
rect 203966 14714 203994 100044
rect 203966 14681 203994 14686
rect 204526 3794 204554 100044
rect 205086 21434 205114 100044
rect 205086 21401 205114 21406
rect 205646 6314 205674 100044
rect 205646 6281 205674 6286
rect 206206 3850 206234 100044
rect 206766 17234 206794 100044
rect 207326 76034 207354 100044
rect 207326 76001 207354 76006
rect 206766 17201 206794 17206
rect 207046 21434 207074 21439
rect 206206 3817 206234 3822
rect 204526 3761 204554 3766
rect 204750 3794 204778 3799
rect 203742 2081 203770 2086
rect 204750 240 204778 3766
rect 206598 3066 206626 3071
rect 205702 2114 205730 2119
rect 205702 240 205730 2086
rect 206598 240 206626 3038
rect 207046 2114 207074 21406
rect 207886 18074 207914 100044
rect 207886 18041 207914 18046
rect 207942 98826 207970 98831
rect 207942 8050 207970 98798
rect 208446 28154 208474 100044
rect 208446 28121 208474 28126
rect 209006 15610 209034 100044
rect 209006 15577 209034 15582
rect 207942 8017 207970 8022
rect 207046 2081 207074 2086
rect 207494 7994 207522 7999
rect 207494 240 207522 7966
rect 209566 7266 209594 100044
rect 210126 29834 210154 100044
rect 210126 29801 210154 29806
rect 209566 7233 209594 7238
rect 210350 9730 210378 9735
rect 209510 3850 209538 3855
rect 208558 2114 208586 2119
rect 208558 240 208586 2086
rect 209510 240 209538 3822
rect 203686 196 203812 240
rect 202748 -480 202860 196
rect 203700 -480 203812 196
rect 204652 196 204778 240
rect 205604 196 205730 240
rect 204652 -480 204764 196
rect 205604 -480 205716 196
rect 206556 -480 206668 240
rect 207494 196 207620 240
rect 207508 -480 207620 196
rect 208460 196 208586 240
rect 209412 196 209538 240
rect 210350 240 210378 9702
rect 210686 8106 210714 100044
rect 211246 8890 211274 100044
rect 211806 22274 211834 100044
rect 212366 98714 212394 100044
rect 212366 98681 212394 98686
rect 211806 22241 211834 22246
rect 212926 9674 212954 100044
rect 213486 14770 213514 100044
rect 214046 98770 214074 100044
rect 214046 98737 214074 98742
rect 213486 14737 213514 14742
rect 212926 9641 212954 9646
rect 213206 12250 213234 12255
rect 211246 8857 211274 8862
rect 210686 8073 210714 8078
rect 212254 6314 212282 6319
rect 211414 2170 211442 2175
rect 211414 240 211442 2142
rect 210350 196 210476 240
rect 208460 -480 208572 196
rect 209412 -480 209524 196
rect 210364 -480 210476 196
rect 211316 196 211442 240
rect 212254 240 212282 6286
rect 213206 240 213234 12222
rect 214606 6370 214634 100044
rect 214662 98770 214690 98775
rect 214662 12194 214690 98742
rect 215166 23954 215194 100044
rect 215166 23921 215194 23926
rect 214662 12161 214690 12166
rect 214606 6337 214634 6342
rect 215222 2954 215250 2959
rect 214270 2226 214298 2231
rect 214270 240 214298 2198
rect 215222 240 215250 2926
rect 215726 2842 215754 100044
rect 216286 98826 216314 100044
rect 216286 98793 216314 98798
rect 216398 99106 216426 99111
rect 216286 98714 216314 98719
rect 215726 2809 215754 2814
rect 216174 4634 216202 4639
rect 216174 240 216202 4606
rect 216286 2954 216314 98686
rect 216398 18914 216426 99078
rect 216846 24794 216874 100044
rect 216846 24761 216874 24766
rect 216398 18881 216426 18886
rect 216286 2921 216314 2926
rect 217406 2898 217434 100044
rect 217966 99106 217994 100044
rect 217966 99073 217994 99078
rect 218526 25634 218554 100044
rect 218526 25601 218554 25606
rect 219086 7154 219114 100044
rect 219646 98770 219674 100044
rect 219646 98737 219674 98742
rect 220206 10514 220234 100044
rect 220766 42434 220794 100044
rect 220766 42401 220794 42406
rect 221326 13034 221354 100044
rect 221326 13001 221354 13006
rect 221382 98322 221410 98327
rect 220206 10481 220234 10486
rect 219086 7121 219114 7126
rect 220822 7154 220850 7159
rect 218918 6370 218946 6375
rect 217406 2865 217434 2870
rect 218078 2954 218106 2959
rect 217126 2282 217154 2287
rect 217126 240 217154 2254
rect 218078 240 218106 2926
rect 212254 196 212380 240
rect 213206 196 213332 240
rect 211316 -480 211428 196
rect 212268 -480 212380 196
rect 213220 -480 213332 196
rect 214172 196 214298 240
rect 215124 196 215250 240
rect 216076 196 216202 240
rect 217028 196 217154 240
rect 217980 196 218106 240
rect 218918 240 218946 6342
rect 219982 2338 220010 2343
rect 219982 240 220010 2310
rect 218918 196 219044 240
rect 214172 -480 214284 196
rect 215124 -480 215236 196
rect 216076 -480 216188 196
rect 217028 -480 217140 196
rect 217980 -480 218092 196
rect 218932 -480 219044 196
rect 219884 196 220010 240
rect 220822 240 220850 7126
rect 221382 3794 221410 98294
rect 221886 16394 221914 100044
rect 221886 16361 221914 16366
rect 222446 8834 222474 100044
rect 222446 8801 222474 8806
rect 222726 98770 222754 98775
rect 221382 3761 221410 3766
rect 221886 3010 221914 3015
rect 221886 240 221914 2982
rect 220822 196 220948 240
rect 219884 -480 219996 196
rect 220836 -480 220948 196
rect 221788 196 221914 240
rect 222726 240 222754 98742
rect 223006 98322 223034 100044
rect 223006 98289 223034 98294
rect 223566 21434 223594 100044
rect 223566 21401 223594 21406
rect 223790 3794 223818 3799
rect 223790 240 223818 3766
rect 224126 3066 224154 100044
rect 224126 3033 224154 3038
rect 224630 97034 224658 97039
rect 222726 196 222852 240
rect 221788 -480 221900 196
rect 222740 -480 222852 196
rect 223692 196 223818 240
rect 224630 240 224658 97006
rect 224686 7994 224714 100044
rect 224686 7961 224714 7966
rect 225246 2114 225274 100044
rect 225806 3850 225834 100044
rect 226366 9730 226394 100044
rect 226366 9697 226394 9702
rect 226534 97874 226562 97879
rect 225806 3817 225834 3822
rect 225246 2081 225274 2086
rect 225694 2114 225722 2119
rect 225694 240 225722 2086
rect 224630 196 224756 240
rect 223692 -480 223804 196
rect 224644 -480 224756 196
rect 225596 196 225722 240
rect 226534 240 226562 97846
rect 226926 2170 226954 100044
rect 227486 6314 227514 100044
rect 228046 12250 228074 100044
rect 228046 12217 228074 12222
rect 228102 99106 228130 99111
rect 227486 6281 227514 6286
rect 228102 3010 228130 99078
rect 228102 2977 228130 2982
rect 228494 98826 228522 98831
rect 226926 2137 226954 2142
rect 227598 2170 227626 2175
rect 227598 240 227626 2142
rect 228494 240 228522 98798
rect 228606 2226 228634 100044
rect 229166 98714 229194 100044
rect 229166 98681 229194 98686
rect 229726 4634 229754 100044
rect 229726 4601 229754 4606
rect 228606 2193 228634 2198
rect 229502 3010 229530 3015
rect 229502 240 229530 2982
rect 230286 2282 230314 100044
rect 230846 2954 230874 100044
rect 231406 6370 231434 100044
rect 231406 6337 231434 6342
rect 230846 2921 230874 2926
rect 231966 2338 231994 100044
rect 232526 7154 232554 100044
rect 233086 99106 233114 100044
rect 233086 99073 233114 99078
rect 233534 99106 233562 99111
rect 233534 97034 233562 99078
rect 233646 98770 233674 100044
rect 233646 98737 233674 98742
rect 233534 97001 233562 97006
rect 234150 98714 234178 98719
rect 232526 7121 232554 7126
rect 231966 2305 231994 2310
rect 232246 6314 232274 6319
rect 230286 2249 230314 2254
rect 231406 2282 231434 2287
rect 230454 2226 230482 2231
rect 230454 240 230482 2198
rect 231406 240 231434 2254
rect 226534 196 226660 240
rect 225596 -480 225708 196
rect 226548 -480 226660 196
rect 227500 196 227626 240
rect 227500 -480 227612 196
rect 228452 -480 228564 240
rect 229404 196 229530 240
rect 230356 196 230482 240
rect 231308 196 231434 240
rect 232246 240 232274 6286
rect 233310 2338 233338 2343
rect 233310 240 233338 2310
rect 232246 196 232372 240
rect 229404 -480 229516 196
rect 230356 -480 230468 196
rect 231308 -480 231420 196
rect 232260 -480 232372 196
rect 233212 196 233338 240
rect 234150 240 234178 98686
rect 234206 3794 234234 100044
rect 234766 99106 234794 100044
rect 234766 99073 234794 99078
rect 234206 3761 234234 3766
rect 235158 2954 235186 2959
rect 235158 240 235186 2926
rect 235326 2114 235354 100044
rect 235886 97874 235914 100044
rect 235886 97841 235914 97846
rect 236446 2170 236474 100044
rect 237006 98826 237034 100044
rect 237006 98793 237034 98798
rect 237566 3010 237594 100044
rect 237566 2977 237594 2982
rect 238070 2394 238098 2399
rect 236446 2137 236474 2142
rect 237118 2170 237146 2175
rect 235326 2081 235354 2086
rect 236166 2114 236194 2119
rect 236166 240 236194 2086
rect 237118 240 237146 2142
rect 238070 240 238098 2366
rect 238126 2226 238154 100044
rect 238686 2282 238714 100044
rect 239246 6314 239274 100044
rect 239246 6281 239274 6286
rect 239806 2338 239834 100044
rect 239806 2305 239834 2310
rect 239862 99050 239890 99055
rect 238686 2249 238714 2254
rect 238126 2193 238154 2198
rect 239022 2226 239050 2231
rect 239022 240 239050 2198
rect 234150 196 234276 240
rect 233212 -480 233324 196
rect 234164 -480 234276 196
rect 235116 -480 235228 240
rect 236068 196 236194 240
rect 237020 196 237146 240
rect 237972 196 238098 240
rect 238924 196 239050 240
rect 239862 240 239890 99022
rect 240366 98714 240394 100044
rect 240366 98681 240394 98686
rect 240814 99106 240842 99111
rect 240814 240 240842 99078
rect 240926 2954 240954 100044
rect 240926 2921 240954 2926
rect 241486 2114 241514 100044
rect 242046 2170 242074 100044
rect 242606 2394 242634 100044
rect 242606 2361 242634 2366
rect 242830 2506 242858 2511
rect 242046 2137 242074 2142
rect 241486 2081 241514 2086
rect 241878 2114 241906 2119
rect 241878 240 241906 2086
rect 242830 240 242858 2478
rect 243166 2226 243194 100044
rect 243726 99050 243754 100044
rect 244286 99106 244314 100044
rect 244286 99073 244314 99078
rect 243726 99017 243754 99022
rect 243166 2193 243194 2198
rect 243670 98378 243698 98383
rect 239862 196 239988 240
rect 240814 196 240940 240
rect 236068 -480 236180 196
rect 237020 -480 237132 196
rect 237972 -480 238084 196
rect 238924 -480 239036 196
rect 239876 -480 239988 196
rect 240828 -480 240940 196
rect 241780 196 241906 240
rect 242732 196 242858 240
rect 243670 240 243698 98350
rect 244622 98322 244650 98327
rect 244622 240 244650 98294
rect 244846 2114 244874 100044
rect 245406 2506 245434 100044
rect 245406 2473 245434 2478
rect 245574 99106 245602 99111
rect 244846 2081 244874 2086
rect 245574 240 245602 99078
rect 245966 98378 245994 100044
rect 245966 98345 245994 98350
rect 246526 98322 246554 100044
rect 247086 99106 247114 100044
rect 247086 99073 247114 99078
rect 247478 99106 247506 99111
rect 246526 98289 246554 98294
rect 246582 99050 246610 99055
rect 246582 240 246610 99022
rect 247478 240 247506 99078
rect 247646 99050 247674 100044
rect 248206 99106 248234 100044
rect 248206 99073 248234 99078
rect 248654 100030 248780 100058
rect 247646 99017 247674 99022
rect 248654 98294 248682 100030
rect 248430 98266 248682 98294
rect 248430 240 248458 98266
rect 249326 10094 249354 100044
rect 249326 10066 249410 10094
rect 249382 240 249410 10066
rect 249886 2114 249914 100044
rect 250446 98322 250474 100044
rect 251006 98378 251034 100044
rect 251566 99106 251594 100044
rect 251566 99073 251594 99078
rect 252126 99050 252154 100044
rect 252126 99017 252154 99022
rect 251006 98345 251034 98350
rect 252238 98378 252266 98383
rect 250446 98289 250474 98294
rect 251286 98322 251314 98327
rect 249886 2081 249914 2086
rect 250334 2114 250362 2119
rect 250334 240 250362 2086
rect 251286 240 251314 98294
rect 252238 240 252266 98350
rect 252686 2170 252714 100044
rect 252686 2137 252714 2142
rect 253190 99106 253218 99111
rect 253190 240 253218 99078
rect 253246 98994 253274 100044
rect 253246 98961 253274 98966
rect 253806 98434 253834 100044
rect 253806 98401 253834 98406
rect 254142 99050 254170 99055
rect 254142 240 254170 99022
rect 254366 2506 254394 100044
rect 254366 2473 254394 2478
rect 254926 2114 254954 100044
rect 255486 98770 255514 100044
rect 256046 99106 256074 100044
rect 256046 99073 256074 99078
rect 255486 98737 255514 98742
rect 255990 98994 256018 98999
rect 255990 92414 256018 98966
rect 256606 98714 256634 100044
rect 256606 98681 256634 98686
rect 256662 99106 256690 99111
rect 255990 92386 256074 92414
rect 254926 2081 254954 2086
rect 255094 2170 255122 2175
rect 255094 240 255122 2142
rect 256046 240 256074 92386
rect 256662 2954 256690 99078
rect 256662 2921 256690 2926
rect 257054 98434 257082 98439
rect 257054 240 257082 98406
rect 257166 2058 257194 100044
rect 257726 99106 257754 100044
rect 257726 99073 257754 99078
rect 258286 51674 258314 100044
rect 258286 51641 258314 51646
rect 258342 99106 258370 99111
rect 258342 3906 258370 99078
rect 258342 3873 258370 3878
rect 257166 2025 257194 2030
rect 257950 2506 257978 2511
rect 257950 240 257978 2478
rect 258846 2170 258874 100044
rect 259406 6314 259434 100044
rect 259406 6281 259434 6286
rect 259854 98770 259882 98775
rect 258846 2137 258874 2142
rect 258902 2114 258930 2119
rect 258902 240 258930 2086
rect 259854 240 259882 98742
rect 259966 7154 259994 100044
rect 259966 7121 259994 7126
rect 260526 2114 260554 100044
rect 261086 3010 261114 100044
rect 261646 99106 261674 100044
rect 261646 99073 261674 99078
rect 261086 2977 261114 2982
rect 261758 98714 261786 98719
rect 260526 2081 260554 2086
rect 260806 2954 260834 2959
rect 260806 240 260834 2926
rect 261758 240 261786 98686
rect 262206 21434 262234 100044
rect 262206 21401 262234 21406
rect 262486 99106 262514 99111
rect 262486 3850 262514 99078
rect 262766 98826 262794 100044
rect 262766 98793 262794 98798
rect 262486 3817 262514 3822
rect 263326 3794 263354 100044
rect 263886 99050 263914 100044
rect 264446 99106 264474 100044
rect 264446 99073 264474 99078
rect 263886 99017 263914 99022
rect 264614 51674 264642 51679
rect 263326 3761 263354 3766
rect 263662 3906 263690 3911
rect 262710 2058 262738 2063
rect 262710 240 262738 2030
rect 263662 240 263690 3878
rect 264614 240 264642 51646
rect 265006 7994 265034 100044
rect 265398 99106 265426 99111
rect 265062 99050 265090 99055
rect 265062 51674 265090 99022
rect 265398 97930 265426 99078
rect 265566 99106 265594 100044
rect 265566 99073 265594 99078
rect 266126 98714 266154 100044
rect 266126 98681 266154 98686
rect 265398 97897 265426 97902
rect 265062 51641 265090 51646
rect 265006 7961 265034 7966
rect 266518 6314 266546 6319
rect 265566 2170 265594 2175
rect 265566 240 265594 2142
rect 266518 240 266546 6286
rect 266686 2954 266714 100044
rect 266742 99106 266770 99111
rect 266742 93674 266770 99078
rect 266742 93641 266770 93646
rect 267246 27314 267274 100044
rect 267806 98770 267834 100044
rect 267806 98737 267834 98742
rect 267246 27281 267274 27286
rect 266686 2921 266714 2926
rect 267470 7154 267498 7159
rect 267470 240 267498 7126
rect 268366 6314 268394 100044
rect 268926 44114 268954 100044
rect 269486 97034 269514 100044
rect 269486 97001 269514 97006
rect 270046 96194 270074 100044
rect 270046 96161 270074 96166
rect 270102 98826 270130 98831
rect 268926 44081 268954 44086
rect 268366 6281 268394 6286
rect 269374 3010 269402 3015
rect 268422 2114 268450 2119
rect 268422 240 268450 2086
rect 269374 240 269402 2982
rect 270102 2562 270130 98798
rect 270102 2529 270130 2534
rect 270326 3850 270354 3855
rect 270326 240 270354 3822
rect 270606 2338 270634 100044
rect 271166 97874 271194 100044
rect 271166 97841 271194 97846
rect 270606 2305 270634 2310
rect 271334 21434 271362 21439
rect 271334 240 271362 21406
rect 271726 7154 271754 100044
rect 271726 7121 271754 7126
rect 272230 2562 272258 2567
rect 272230 240 272258 2534
rect 272286 2282 272314 100044
rect 272286 2249 272314 2254
rect 272846 2226 272874 100044
rect 272846 2193 272874 2198
rect 273182 3794 273210 3799
rect 273182 240 273210 3766
rect 273406 2170 273434 100044
rect 273406 2137 273434 2142
rect 273966 2114 273994 100044
rect 275926 98770 275954 98775
rect 275086 97930 275114 97935
rect 273966 2081 273994 2086
rect 274134 51674 274162 51679
rect 274134 240 274162 51646
rect 275086 240 275114 97902
rect 275926 3010 275954 98742
rect 277942 98714 277970 98719
rect 276990 93674 277018 93679
rect 275926 2977 275954 2982
rect 276038 7994 276066 7999
rect 276038 240 276066 7966
rect 276990 240 277018 93646
rect 277942 240 277970 98686
rect 282198 82866 282226 104902
rect 286510 97874 286538 97879
rect 282198 82833 282226 82838
rect 283654 97034 283682 97039
rect 282702 44114 282730 44119
rect 279846 27314 279874 27319
rect 278894 2954 278922 2959
rect 278894 240 278922 2926
rect 279846 240 279874 27286
rect 281750 6314 281778 6319
rect 280798 3010 280826 3015
rect 280798 240 280826 2982
rect 281750 240 281778 6286
rect 282702 240 282730 44086
rect 283654 240 283682 97006
rect 284606 96194 284634 96199
rect 284606 240 284634 96166
rect 285614 2338 285642 2343
rect 285614 240 285642 2310
rect 286510 240 286538 97846
rect 287462 7154 287490 7159
rect 287462 240 287490 7126
rect 288414 2282 288442 2287
rect 288414 240 288442 2254
rect 290318 2226 290346 2231
rect 290318 240 290346 2198
rect 291270 2170 291298 2175
rect 291270 240 291298 2142
rect 292222 2114 292250 2119
rect 292222 240 292250 2086
rect 243670 196 243796 240
rect 244622 196 244748 240
rect 245574 196 245700 240
rect 241780 -480 241892 196
rect 242732 -480 242844 196
rect 243684 -480 243796 196
rect 244636 -480 244748 196
rect 245588 -480 245700 196
rect 246540 -480 246652 240
rect 247478 196 247604 240
rect 248430 196 248556 240
rect 249382 196 249508 240
rect 250334 196 250460 240
rect 251286 196 251412 240
rect 252238 196 252364 240
rect 253190 196 253316 240
rect 254142 196 254268 240
rect 255094 196 255220 240
rect 256046 196 256172 240
rect 247492 -480 247604 196
rect 248444 -480 248556 196
rect 249396 -480 249508 196
rect 250348 -480 250460 196
rect 251300 -480 251412 196
rect 252252 -480 252364 196
rect 253204 -480 253316 196
rect 254156 -480 254268 196
rect 255108 -480 255220 196
rect 256060 -480 256172 196
rect 257012 -480 257124 240
rect 257950 196 258076 240
rect 258902 196 259028 240
rect 259854 196 259980 240
rect 260806 196 260932 240
rect 261758 196 261884 240
rect 262710 196 262836 240
rect 263662 196 263788 240
rect 264614 196 264740 240
rect 265566 196 265692 240
rect 266518 196 266644 240
rect 267470 196 267596 240
rect 268422 196 268548 240
rect 269374 196 269500 240
rect 270326 196 270452 240
rect 257964 -480 258076 196
rect 258916 -480 259028 196
rect 259868 -480 259980 196
rect 260820 -480 260932 196
rect 261772 -480 261884 196
rect 262724 -480 262836 196
rect 263676 -480 263788 196
rect 264628 -480 264740 196
rect 265580 -480 265692 196
rect 266532 -480 266644 196
rect 267484 -480 267596 196
rect 268436 -480 268548 196
rect 269388 -480 269500 196
rect 270340 -480 270452 196
rect 271292 -480 271404 240
rect 272230 196 272356 240
rect 273182 196 273308 240
rect 274134 196 274260 240
rect 275086 196 275212 240
rect 276038 196 276164 240
rect 276990 196 277116 240
rect 277942 196 278068 240
rect 278894 196 279020 240
rect 279846 196 279972 240
rect 280798 196 280924 240
rect 281750 196 281876 240
rect 282702 196 282828 240
rect 283654 196 283780 240
rect 284606 196 284732 240
rect 272244 -480 272356 196
rect 273196 -480 273308 196
rect 274148 -480 274260 196
rect 275100 -480 275212 196
rect 276052 -480 276164 196
rect 277004 -480 277116 196
rect 277956 -480 278068 196
rect 278908 -480 279020 196
rect 279860 -480 279972 196
rect 280812 -480 280924 196
rect 281764 -480 281876 196
rect 282716 -480 282828 196
rect 283668 -480 283780 196
rect 284620 -480 284732 196
rect 285572 -480 285684 240
rect 286510 196 286636 240
rect 287462 196 287588 240
rect 288414 196 288540 240
rect 286524 -480 286636 196
rect 287476 -480 287588 196
rect 288428 -480 288540 196
rect 289380 -480 289492 240
rect 290318 196 290444 240
rect 291270 196 291396 240
rect 292222 196 292348 240
rect 290332 -480 290444 196
rect 291284 -480 291396 196
rect 292236 -480 292348 196
<< via2 >>
rect 98686 238014 98714 238042
rect 281414 156310 281442 156338
rect 281414 155526 281442 155554
rect 98686 131278 98714 131306
rect 281470 126854 281498 126882
rect 281470 122486 281498 122514
rect 282142 119294 282170 119322
rect 282142 102662 282170 102690
rect 282198 104902 282226 104930
rect 104566 98910 104594 98938
rect 96166 98798 96194 98826
rect 58366 98742 58394 98770
rect 5670 98686 5698 98714
rect 11382 97846 11410 97874
rect 6622 27286 6650 27314
rect 7574 9646 7602 9674
rect 8638 3766 8666 3794
rect 10542 2142 10570 2170
rect 9590 2086 9618 2114
rect 15190 97006 15218 97034
rect 14294 61726 14322 61754
rect 13398 4606 13426 4634
rect 12446 3822 12474 3850
rect 43750 96166 43778 96194
rect 24710 86926 24738 86954
rect 17094 84406 17122 84434
rect 16254 4662 16282 4690
rect 21406 81046 21434 81074
rect 18998 54166 19026 54194
rect 18158 2198 18186 2226
rect 20902 14686 20930 14714
rect 20062 2030 20090 2058
rect 22806 80206 22834 80234
rect 21406 2030 21434 2058
rect 21966 2254 21994 2282
rect 23758 52486 23786 52514
rect 26614 79366 26642 79394
rect 25774 2310 25802 2338
rect 29470 78526 29498 78554
rect 28574 28126 28602 28154
rect 27566 26446 27594 26474
rect 32326 77686 32354 77714
rect 31374 42406 31402 42434
rect 30422 33166 30450 33194
rect 35182 76006 35210 76034
rect 34230 15526 34258 15554
rect 33390 5446 33418 5474
rect 38038 75166 38066 75194
rect 37086 48286 37114 48314
rect 36134 6286 36162 6314
rect 39942 66766 39970 66794
rect 38990 6342 39018 6370
rect 42854 64246 42882 64274
rect 41846 7126 41874 7154
rect 41006 3878 41034 3906
rect 46606 93646 46634 93674
rect 44702 34006 44730 34034
rect 45654 7182 45682 7210
rect 52318 92806 52346 92834
rect 51366 58366 51394 58394
rect 47558 55006 47586 55034
rect 48510 43246 48538 43274
rect 50414 13006 50442 13034
rect 49518 2982 49546 3010
rect 55174 91126 55202 91154
rect 53270 34846 53298 34874
rect 54222 7966 54250 7994
rect 56126 56686 56154 56714
rect 57134 8022 57162 8050
rect 86590 97902 86618 97930
rect 68502 97062 68530 97090
rect 66598 90286 66626 90314
rect 64694 72646 64722 72674
rect 62790 70126 62818 70154
rect 61838 44926 61866 44954
rect 58366 2982 58394 3010
rect 58982 30646 59010 30674
rect 58142 2926 58170 2954
rect 59934 8078 59962 8106
rect 60998 2982 61026 3010
rect 63798 3038 63826 3066
rect 65646 12166 65674 12194
rect 67550 57526 67578 57554
rect 69454 89446 69482 89474
rect 72310 87766 72338 87794
rect 71414 8806 71442 8834
rect 70406 6398 70434 6426
rect 75166 86982 75194 87010
rect 73262 71806 73290 71834
rect 74214 8862 74242 8890
rect 78022 85246 78050 85274
rect 76118 70966 76146 70994
rect 77070 37366 77098 37394
rect 83734 84462 83762 84490
rect 82782 53326 82810 53354
rect 81830 18886 81858 18914
rect 80878 12222 80906 12250
rect 78974 9702 79002 9730
rect 79926 8918 79954 8946
rect 85694 44086 85722 44114
rect 84686 7238 84714 7266
rect 91350 92862 91378 92890
rect 89446 88606 89474 88634
rect 87542 65926 87570 65954
rect 88494 60046 88522 60074
rect 90398 36526 90426 36554
rect 94206 91182 94234 91210
rect 92302 81102 92330 81130
rect 93254 51646 93282 51674
rect 96110 22246 96138 22274
rect 95270 2534 95298 2562
rect 96166 2534 96194 2562
rect 98014 96222 98042 96250
rect 97174 1246 97202 1274
rect 103726 93702 103754 93730
rect 100870 81886 100898 81914
rect 99974 39046 100002 39074
rect 98966 18046 98994 18074
rect 101822 69286 101850 69314
rect 102774 39886 102802 39914
rect 105798 98854 105826 98882
rect 104566 12222 104594 12250
rect 104678 35686 104706 35714
rect 105630 21406 105658 21434
rect 105966 98686 105994 98714
rect 106526 27286 106554 27314
rect 107086 9646 107114 9674
rect 107534 9646 107562 9674
rect 105798 2534 105826 2562
rect 106582 2534 106610 2562
rect 107646 3766 107674 3794
rect 108206 2086 108234 2114
rect 108486 29806 108514 29834
rect 109326 97846 109354 97874
rect 108766 2142 108794 2170
rect 109438 13062 109466 13090
rect 111566 97006 111594 97034
rect 111006 61726 111034 61754
rect 111342 24766 111370 24794
rect 110446 4606 110474 4634
rect 110502 4718 110530 4746
rect 109886 3822 109914 3850
rect 112686 84406 112714 84434
rect 112126 4662 112154 4690
rect 112406 3766 112434 3794
rect 114366 81046 114394 81074
rect 113806 54166 113834 54194
rect 114254 23926 114282 23954
rect 113246 2198 113274 2226
rect 113302 16366 113330 16394
rect 114926 14686 114954 14714
rect 115150 14686 115178 14714
rect 116046 80206 116074 80234
rect 116606 52486 116634 52514
rect 117054 97006 117082 97034
rect 115486 2254 115514 2282
rect 116102 25606 116130 25634
rect 117166 86926 117194 86954
rect 118286 79366 118314 79394
rect 119966 78526 119994 78554
rect 121646 77686 121674 77714
rect 121086 42406 121114 42434
rect 120526 33166 120554 33194
rect 119406 28126 119434 28154
rect 121814 27286 121842 27314
rect 118846 26446 118874 26474
rect 118958 26446 118986 26474
rect 117726 2310 117754 2338
rect 118006 12222 118034 12250
rect 119910 17262 119938 17290
rect 120862 15582 120890 15610
rect 123326 76006 123354 76034
rect 122766 15526 122794 15554
rect 123718 17206 123746 17234
rect 122206 5446 122234 5474
rect 122878 3822 122906 3850
rect 124278 98294 124306 98322
rect 124278 96166 124306 96194
rect 125006 75166 125034 75194
rect 124446 48286 124474 48314
rect 123886 6286 123914 6314
rect 124670 10486 124698 10514
rect 126126 66766 126154 66794
rect 125566 6342 125594 6370
rect 126574 18102 126602 18130
rect 125734 4606 125762 4634
rect 128366 98294 128394 98322
rect 127806 64246 127834 64274
rect 127246 7126 127274 7154
rect 128534 34062 128562 34090
rect 126686 3878 126714 3906
rect 127526 6286 127554 6314
rect 128926 34006 128954 34034
rect 129430 18942 129458 18970
rect 130046 93646 130074 93674
rect 130606 55006 130634 55034
rect 131726 98742 131754 98770
rect 131166 43246 131194 43274
rect 129486 7182 129514 7210
rect 130382 28126 130410 28154
rect 131334 16422 131362 16450
rect 133406 92806 133434 92834
rect 132846 58366 132874 58394
rect 133966 34846 133994 34874
rect 134190 33166 134218 33194
rect 132286 13006 132314 13034
rect 132342 21462 132370 21490
rect 133238 15526 133266 15554
rect 135086 91126 135114 91154
rect 135646 56686 135674 56714
rect 135702 98686 135730 98714
rect 135702 12166 135730 12194
rect 136206 8022 136234 8050
rect 134526 7966 134554 7994
rect 136094 7126 136122 7154
rect 135198 3878 135226 3906
rect 136766 2926 136794 2954
rect 137046 30702 137074 30730
rect 137382 98294 137410 98322
rect 137382 72646 137410 72674
rect 137326 30646 137354 30674
rect 137886 8078 137914 8106
rect 137998 7966 138026 7994
rect 139062 98966 139090 98994
rect 139062 90286 139090 90314
rect 139566 70126 139594 70154
rect 139006 44926 139034 44954
rect 138446 2982 138474 3010
rect 138950 22302 138978 22330
rect 140014 5446 140042 5474
rect 141806 98966 141834 98994
rect 141246 98686 141274 98714
rect 140686 98294 140714 98322
rect 142422 99078 142450 99106
rect 143486 99078 143514 99106
rect 142758 97062 142786 97090
rect 142422 89446 142450 89474
rect 142366 57526 142394 57554
rect 143710 64246 143738 64274
rect 140126 3038 140154 3066
rect 141918 3038 141946 3066
rect 140966 2926 140994 2954
rect 142870 2982 142898 3010
rect 145166 87766 145194 87794
rect 145670 71806 145698 71834
rect 145726 98686 145754 98714
rect 145614 13006 145642 13034
rect 144606 8806 144634 8834
rect 144662 8974 144690 9002
rect 144046 6398 144074 6426
rect 146846 86982 146874 87010
rect 147406 70966 147434 70994
rect 147518 97846 147546 97874
rect 146286 8862 146314 8890
rect 145726 2982 145754 3010
rect 146566 6342 146594 6370
rect 148526 85246 148554 85274
rect 147966 37366 147994 37394
rect 148470 14742 148498 14770
rect 149086 9702 149114 9730
rect 149422 9702 149450 9730
rect 150206 98910 150234 98938
rect 149646 8918 149674 8946
rect 150374 23982 150402 24010
rect 151886 84462 151914 84490
rect 151326 53326 151354 53354
rect 150766 18886 150794 18914
rect 151326 18886 151354 18914
rect 153566 97902 153594 97930
rect 154182 99022 154210 99050
rect 154182 92862 154210 92890
rect 154126 65926 154154 65954
rect 154182 65982 154210 66010
rect 153006 44086 153034 44114
rect 152446 7238 152474 7266
rect 153230 8022 153258 8050
rect 152278 7182 152306 7210
rect 155246 88606 155274 88634
rect 154686 60046 154714 60074
rect 155862 99078 155890 99106
rect 156926 99078 156954 99106
rect 156366 99022 156394 99050
rect 155862 81102 155890 81130
rect 157486 51646 157514 51674
rect 157542 99078 157570 99106
rect 155806 36526 155834 36554
rect 157094 25662 157122 25690
rect 156086 24822 156114 24850
rect 155134 8806 155162 8834
rect 159166 99078 159194 99106
rect 158606 98798 158634 98826
rect 159166 98742 159194 98770
rect 157654 91182 157682 91210
rect 157542 22246 157570 22274
rect 158942 6398 158970 6426
rect 158102 2534 158130 2562
rect 159166 2534 159194 2562
rect 160286 96222 160314 96250
rect 161966 81886 161994 81914
rect 162526 69286 162554 69314
rect 162750 69286 162778 69314
rect 161406 39046 161434 39074
rect 160846 18046 160874 18074
rect 160846 12166 160874 12194
rect 159726 1246 159754 1274
rect 159894 10542 159922 10570
rect 161798 9758 161826 9786
rect 163646 93702 163674 93730
rect 163086 39886 163114 39914
rect 164206 35686 164234 35714
rect 165326 98854 165354 98882
rect 164766 21406 164794 21434
rect 165606 12278 165634 12306
rect 164766 4662 164794 4690
rect 163758 3038 163786 3066
rect 165886 9646 165914 9674
rect 165942 98798 165970 98826
rect 166446 29806 166474 29834
rect 165942 3878 165970 3906
rect 166558 13118 166586 13146
rect 167006 13062 167034 13090
rect 168126 24766 168154 24794
rect 168462 26502 168490 26530
rect 167566 4718 167594 4746
rect 167622 3878 167650 3906
rect 169302 99022 169330 99050
rect 169806 23926 169834 23954
rect 169302 17262 169330 17290
rect 169246 16366 169274 16394
rect 169414 16366 169442 16394
rect 168686 3766 168714 3794
rect 170926 25606 170954 25634
rect 170982 99078 171010 99106
rect 170366 14686 170394 14714
rect 170422 17262 170450 17290
rect 172046 99078 172074 99106
rect 171318 97006 171346 97034
rect 172606 26446 172634 26474
rect 172662 99078 172690 99106
rect 173726 99078 173754 99106
rect 173166 99022 173194 99050
rect 172662 15582 172690 15610
rect 172718 27342 172746 27370
rect 170982 12222 171010 12250
rect 172270 14686 172298 14714
rect 171430 2086 171458 2114
rect 174286 27286 174314 27314
rect 174342 98966 174370 98994
rect 174174 21406 174202 21434
rect 172718 2086 172746 2114
rect 173334 3766 173362 3794
rect 174342 6286 174370 6314
rect 175406 17206 175434 17234
rect 175966 10486 175994 10514
rect 176022 99078 176050 99106
rect 174846 3822 174874 3850
rect 175126 6286 175154 6314
rect 176526 99078 176554 99106
rect 177646 98966 177674 98994
rect 177646 98854 177674 98882
rect 177646 30702 177674 30730
rect 177982 76006 178010 76034
rect 177086 18102 177114 18130
rect 176022 4606 176050 4634
rect 177030 17206 177058 17234
rect 176190 3822 176218 3850
rect 178206 34062 178234 34090
rect 179326 28126 179354 28154
rect 179382 99078 179410 99106
rect 178766 18942 178794 18970
rect 178934 18046 178962 18074
rect 179886 99078 179914 99106
rect 180446 21462 180474 21490
rect 179382 16422 179410 16450
rect 180838 15582 180866 15610
rect 179998 2086 180026 2114
rect 182126 98798 182154 98826
rect 181566 33166 181594 33194
rect 181006 15526 181034 15554
rect 181790 7238 181818 7266
rect 183246 98854 183274 98882
rect 183526 29806 183554 29834
rect 182686 7126 182714 7154
rect 182854 28126 182882 28154
rect 182798 2142 182826 2170
rect 182854 2086 182882 2114
rect 183526 2086 183554 2114
rect 183694 8078 183722 8106
rect 184366 22302 184394 22330
rect 184422 98798 184450 98826
rect 184422 8974 184450 9002
rect 183806 7966 183834 7994
rect 184646 8862 184674 8890
rect 184926 5446 184954 5474
rect 185486 2926 185514 2954
rect 185654 22246 185682 22274
rect 186606 98686 186634 98714
rect 186102 98294 186130 98322
rect 187726 98798 187754 98826
rect 187166 98294 187194 98322
rect 187726 98686 187754 98714
rect 186102 64246 186130 64274
rect 186046 2982 186074 3010
rect 187502 9646 187530 9674
rect 186662 2534 186690 2562
rect 188846 98686 188874 98714
rect 189406 97846 189434 97874
rect 189966 14742 189994 14770
rect 190246 14742 190274 14770
rect 188286 13006 188314 13034
rect 187726 6342 187754 6370
rect 189518 3094 189546 3122
rect 188566 2086 188594 2114
rect 191086 23982 191114 24010
rect 191142 98686 191170 98714
rect 190526 9702 190554 9730
rect 190246 2086 190274 2114
rect 190358 6342 190386 6370
rect 191646 18886 191674 18914
rect 193326 65982 193354 66010
rect 192766 8022 192794 8050
rect 192822 23926 192850 23954
rect 192206 7182 192234 7210
rect 191142 2534 191170 2562
rect 192318 2926 192346 2954
rect 191422 2478 191450 2506
rect 194446 24822 194474 24850
rect 194502 98350 194530 98378
rect 193886 8806 193914 8834
rect 192822 2478 192850 2506
rect 193214 8022 193242 8050
rect 195006 25662 195034 25690
rect 195286 99078 195314 99106
rect 195566 98742 195594 98770
rect 195286 10542 195314 10570
rect 195342 24766 195370 24794
rect 194502 3038 194530 3066
rect 195230 2982 195258 3010
rect 194278 2086 194306 2114
rect 195342 2086 195370 2114
rect 196070 18886 196098 18914
rect 196686 99078 196714 99106
rect 196126 6398 196154 6426
rect 197022 25606 197050 25634
rect 197246 12166 197274 12194
rect 198366 69286 198394 69314
rect 198646 99078 198674 99106
rect 198926 98350 198954 98378
rect 198646 17262 198674 17290
rect 197806 9758 197834 9786
rect 198926 12166 198954 12194
rect 197974 7126 198002 7154
rect 199486 4662 199514 4690
rect 199542 98742 199570 98770
rect 200606 13118 200634 13146
rect 200830 42406 200858 42434
rect 200046 12278 200074 12306
rect 199542 3094 199570 3122
rect 199934 10486 199962 10514
rect 201726 26502 201754 26530
rect 202846 99078 202874 99106
rect 203406 27342 203434 27370
rect 202286 16366 202314 16394
rect 203742 16366 203770 16394
rect 201166 3878 201194 3906
rect 201782 13006 201810 13034
rect 203686 8806 203714 8834
rect 202846 2086 202874 2114
rect 203966 14686 203994 14714
rect 205086 21406 205114 21434
rect 205646 6286 205674 6314
rect 207326 76006 207354 76034
rect 206766 17206 206794 17234
rect 207046 21406 207074 21434
rect 206206 3822 206234 3850
rect 204526 3766 204554 3794
rect 204750 3766 204778 3794
rect 203742 2086 203770 2114
rect 206598 3038 206626 3066
rect 205702 2086 205730 2114
rect 207886 18046 207914 18074
rect 207942 98798 207970 98826
rect 208446 28126 208474 28154
rect 209006 15582 209034 15610
rect 207942 8022 207970 8050
rect 207046 2086 207074 2114
rect 207494 7966 207522 7994
rect 210126 29806 210154 29834
rect 209566 7238 209594 7266
rect 210350 9702 210378 9730
rect 209510 3822 209538 3850
rect 208558 2086 208586 2114
rect 212366 98686 212394 98714
rect 211806 22246 211834 22274
rect 214046 98742 214074 98770
rect 213486 14742 213514 14770
rect 212926 9646 212954 9674
rect 213206 12222 213234 12250
rect 211246 8862 211274 8890
rect 210686 8078 210714 8106
rect 212254 6286 212282 6314
rect 211414 2142 211442 2170
rect 214662 98742 214690 98770
rect 215166 23926 215194 23954
rect 214662 12166 214690 12194
rect 214606 6342 214634 6370
rect 215222 2926 215250 2954
rect 214270 2198 214298 2226
rect 216286 98798 216314 98826
rect 216398 99078 216426 99106
rect 216286 98686 216314 98714
rect 215726 2814 215754 2842
rect 216174 4606 216202 4634
rect 216846 24766 216874 24794
rect 216398 18886 216426 18914
rect 216286 2926 216314 2954
rect 217966 99078 217994 99106
rect 218526 25606 218554 25634
rect 219646 98742 219674 98770
rect 220766 42406 220794 42434
rect 221326 13006 221354 13034
rect 221382 98294 221410 98322
rect 220206 10486 220234 10514
rect 219086 7126 219114 7154
rect 220822 7126 220850 7154
rect 218918 6342 218946 6370
rect 217406 2870 217434 2898
rect 218078 2926 218106 2954
rect 217126 2254 217154 2282
rect 219982 2310 220010 2338
rect 221886 16366 221914 16394
rect 222446 8806 222474 8834
rect 222726 98742 222754 98770
rect 221382 3766 221410 3794
rect 221886 2982 221914 3010
rect 223006 98294 223034 98322
rect 223566 21406 223594 21434
rect 223790 3766 223818 3794
rect 224126 3038 224154 3066
rect 224630 97006 224658 97034
rect 224686 7966 224714 7994
rect 226366 9702 226394 9730
rect 226534 97846 226562 97874
rect 225806 3822 225834 3850
rect 225246 2086 225274 2114
rect 225694 2086 225722 2114
rect 228046 12222 228074 12250
rect 228102 99078 228130 99106
rect 227486 6286 227514 6314
rect 228102 2982 228130 3010
rect 228494 98798 228522 98826
rect 226926 2142 226954 2170
rect 227598 2142 227626 2170
rect 229166 98686 229194 98714
rect 229726 4606 229754 4634
rect 228606 2198 228634 2226
rect 229502 2982 229530 3010
rect 231406 6342 231434 6370
rect 230846 2926 230874 2954
rect 233086 99078 233114 99106
rect 233534 99078 233562 99106
rect 233646 98742 233674 98770
rect 233534 97006 233562 97034
rect 234150 98686 234178 98714
rect 232526 7126 232554 7154
rect 231966 2310 231994 2338
rect 232246 6286 232274 6314
rect 230286 2254 230314 2282
rect 231406 2254 231434 2282
rect 230454 2198 230482 2226
rect 233310 2310 233338 2338
rect 234766 99078 234794 99106
rect 234206 3766 234234 3794
rect 235158 2926 235186 2954
rect 235886 97846 235914 97874
rect 237006 98798 237034 98826
rect 237566 2982 237594 3010
rect 238070 2366 238098 2394
rect 236446 2142 236474 2170
rect 237118 2142 237146 2170
rect 235326 2086 235354 2114
rect 236166 2086 236194 2114
rect 239246 6286 239274 6314
rect 239806 2310 239834 2338
rect 239862 99022 239890 99050
rect 238686 2254 238714 2282
rect 238126 2198 238154 2226
rect 239022 2198 239050 2226
rect 240366 98686 240394 98714
rect 240814 99078 240842 99106
rect 240926 2926 240954 2954
rect 242606 2366 242634 2394
rect 242830 2478 242858 2506
rect 242046 2142 242074 2170
rect 241486 2086 241514 2114
rect 241878 2086 241906 2114
rect 244286 99078 244314 99106
rect 243726 99022 243754 99050
rect 243166 2198 243194 2226
rect 243670 98350 243698 98378
rect 244622 98294 244650 98322
rect 245406 2478 245434 2506
rect 245574 99078 245602 99106
rect 244846 2086 244874 2114
rect 245966 98350 245994 98378
rect 247086 99078 247114 99106
rect 247478 99078 247506 99106
rect 246526 98294 246554 98322
rect 246582 99022 246610 99050
rect 248206 99078 248234 99106
rect 247646 99022 247674 99050
rect 251566 99078 251594 99106
rect 252126 99022 252154 99050
rect 251006 98350 251034 98378
rect 252238 98350 252266 98378
rect 250446 98294 250474 98322
rect 251286 98294 251314 98322
rect 249886 2086 249914 2114
rect 250334 2086 250362 2114
rect 252686 2142 252714 2170
rect 253190 99078 253218 99106
rect 253246 98966 253274 98994
rect 253806 98406 253834 98434
rect 254142 99022 254170 99050
rect 254366 2478 254394 2506
rect 256046 99078 256074 99106
rect 255486 98742 255514 98770
rect 255990 98966 256018 98994
rect 256606 98686 256634 98714
rect 256662 99078 256690 99106
rect 254926 2086 254954 2114
rect 255094 2142 255122 2170
rect 256662 2926 256690 2954
rect 257054 98406 257082 98434
rect 257726 99078 257754 99106
rect 258286 51646 258314 51674
rect 258342 99078 258370 99106
rect 258342 3878 258370 3906
rect 257166 2030 257194 2058
rect 257950 2478 257978 2506
rect 259406 6286 259434 6314
rect 259854 98742 259882 98770
rect 258846 2142 258874 2170
rect 258902 2086 258930 2114
rect 259966 7126 259994 7154
rect 261646 99078 261674 99106
rect 261086 2982 261114 3010
rect 261758 98686 261786 98714
rect 260526 2086 260554 2114
rect 260806 2926 260834 2954
rect 262206 21406 262234 21434
rect 262486 99078 262514 99106
rect 262766 98798 262794 98826
rect 262486 3822 262514 3850
rect 264446 99078 264474 99106
rect 263886 99022 263914 99050
rect 264614 51646 264642 51674
rect 263326 3766 263354 3794
rect 263662 3878 263690 3906
rect 262710 2030 262738 2058
rect 265398 99078 265426 99106
rect 265062 99022 265090 99050
rect 265566 99078 265594 99106
rect 266126 98686 266154 98714
rect 265398 97902 265426 97930
rect 265062 51646 265090 51674
rect 265006 7966 265034 7994
rect 266518 6286 266546 6314
rect 265566 2142 265594 2170
rect 266742 99078 266770 99106
rect 266742 93646 266770 93674
rect 267806 98742 267834 98770
rect 267246 27286 267274 27314
rect 266686 2926 266714 2954
rect 267470 7126 267498 7154
rect 269486 97006 269514 97034
rect 270046 96166 270074 96194
rect 270102 98798 270130 98826
rect 268926 44086 268954 44114
rect 268366 6286 268394 6314
rect 269374 2982 269402 3010
rect 268422 2086 268450 2114
rect 270102 2534 270130 2562
rect 270326 3822 270354 3850
rect 271166 97846 271194 97874
rect 270606 2310 270634 2338
rect 271334 21406 271362 21434
rect 271726 7126 271754 7154
rect 272230 2534 272258 2562
rect 272286 2254 272314 2282
rect 272846 2198 272874 2226
rect 273182 3766 273210 3794
rect 273406 2142 273434 2170
rect 275926 98742 275954 98770
rect 275086 97902 275114 97930
rect 273966 2086 273994 2114
rect 274134 51646 274162 51674
rect 277942 98686 277970 98714
rect 276990 93646 277018 93674
rect 275926 2982 275954 3010
rect 276038 7966 276066 7994
rect 286510 97846 286538 97874
rect 282198 82838 282226 82866
rect 283654 97006 283682 97034
rect 282702 44086 282730 44114
rect 279846 27286 279874 27314
rect 278894 2926 278922 2954
rect 281750 6286 281778 6314
rect 280798 2982 280826 3010
rect 284606 96166 284634 96194
rect 285614 2310 285642 2338
rect 287462 7126 287490 7154
rect 288414 2254 288442 2282
rect 290318 2198 290346 2226
rect 291270 2142 291298 2170
rect 292222 2086 292250 2114
<< metal3 >>
rect 297780 294308 298500 294420
rect -480 293580 240 293692
rect 297780 287700 298500 287812
rect -480 286524 240 286636
rect 297780 281092 298500 281204
rect -480 279468 240 279580
rect 98681 274974 98686 275002
rect 98714 274974 100044 275002
rect 279972 274974 281414 275002
rect 281442 274974 281447 275002
rect 297780 274484 298500 274596
rect -480 272412 240 272524
rect 297780 267876 298500 267988
rect 2081 267582 2086 267610
rect 2114 267582 100044 267610
rect 279972 267582 281806 267610
rect 281834 267582 281839 267610
rect -480 265356 240 265468
rect 297780 261268 298500 261380
rect 98737 260190 98742 260218
rect 98770 260190 100044 260218
rect 279972 260190 281862 260218
rect 281890 260190 281895 260218
rect -480 258300 240 258412
rect 297780 254660 298500 254772
rect 98849 252798 98854 252826
rect 98882 252798 100044 252826
rect 279972 252798 284326 252826
rect 284354 252798 284359 252826
rect -480 251244 240 251356
rect 297780 248052 298500 248164
rect 2137 245406 2142 245434
rect 2170 245406 100044 245434
rect 279972 245406 286846 245434
rect 286874 245406 286879 245434
rect -480 244188 240 244300
rect 297780 241444 298500 241556
rect 98681 238014 98686 238042
rect 98714 238014 100044 238042
rect 279972 238014 281470 238042
rect 281498 238014 281503 238042
rect -480 237132 240 237244
rect 297780 234836 298500 234948
rect 98793 230622 98798 230650
rect 98826 230622 100044 230650
rect 279972 230622 283486 230650
rect 283514 230622 283519 230650
rect -480 230076 240 230188
rect 297780 228228 298500 228340
rect 2193 223230 2198 223258
rect 2226 223230 100044 223258
rect 279972 223230 286006 223258
rect 286034 223230 286039 223258
rect -480 223020 240 223132
rect 297780 221620 298500 221732
rect -480 215964 240 216076
rect 98961 215838 98966 215866
rect 98994 215838 100044 215866
rect 279972 215838 281526 215866
rect 281554 215838 281559 215866
rect 297780 215012 298500 215124
rect -480 208908 240 209020
rect 98905 208446 98910 208474
rect 98938 208446 100044 208474
rect 279972 208446 282646 208474
rect 282674 208446 282679 208474
rect 297780 208404 298500 208516
rect -480 201852 240 201964
rect 297780 201796 298500 201908
rect 3761 201054 3766 201082
rect 3794 201054 100044 201082
rect 279972 201054 292726 201082
rect 292754 201054 292759 201082
rect 297780 195188 298500 195300
rect -480 194796 240 194908
rect 99017 193662 99022 193690
rect 99050 193662 100044 193690
rect 279972 193662 281582 193690
rect 281610 193662 281615 193690
rect 297780 188580 298500 188692
rect -480 187740 240 187852
rect 98625 186270 98630 186298
rect 98658 186270 100044 186298
rect 279972 186270 281918 186298
rect 281946 186270 281951 186298
rect 297780 181972 298500 182084
rect -480 180684 240 180796
rect 2249 178878 2254 178906
rect 2282 178878 100044 178906
rect 279972 178878 289366 178906
rect 289394 178878 289399 178906
rect 297780 175364 298500 175476
rect -480 173628 240 173740
rect 99073 171486 99078 171514
rect 99106 171486 100044 171514
rect 279972 171486 281974 171514
rect 282002 171486 282007 171514
rect 297780 168756 298500 168868
rect -480 166586 240 166684
rect -480 166572 98686 166586
rect 196 166558 98686 166572
rect 98714 166558 98719 166586
rect 98681 164094 98686 164122
rect 98714 164094 100044 164122
rect 279972 164094 282030 164122
rect 282058 164094 282063 164122
rect 297780 162148 298500 162260
rect -480 159586 240 159628
rect -480 159558 2086 159586
rect 2114 159558 2119 159586
rect -480 159516 240 159558
rect 2081 156702 2086 156730
rect 2114 156702 100044 156730
rect 279972 156702 282086 156730
rect 282114 156702 282119 156730
rect 281395 156310 281414 156338
rect 281442 156310 281447 156338
rect 297780 155554 298500 155652
rect 281409 155526 281414 155554
rect 281442 155540 298500 155554
rect 281442 155526 297836 155540
rect -480 152474 240 152572
rect -480 152460 98742 152474
rect 196 152446 98742 152460
rect 98770 152446 98775 152474
rect 98737 149310 98742 149338
rect 98770 149310 100044 149338
rect 279972 149310 282142 149338
rect 282170 149310 282175 149338
rect 297780 148946 298500 149044
rect 281801 148918 281806 148946
rect 281834 148932 298500 148946
rect 281834 148918 297836 148932
rect -480 145418 240 145516
rect -480 145404 98854 145418
rect 196 145390 98854 145404
rect 98882 145390 98887 145418
rect 297780 142338 298500 142436
rect 281857 142310 281862 142338
rect 281890 142324 298500 142338
rect 281890 142310 297836 142324
rect 98849 141918 98854 141946
rect 98882 141918 100044 141946
rect 279972 141918 281806 141946
rect 281834 141918 281839 141946
rect 196 138460 2142 138474
rect -480 138446 2142 138460
rect 2170 138446 2175 138474
rect -480 138348 240 138446
rect 297780 135730 298500 135828
rect 284321 135702 284326 135730
rect 284354 135716 298500 135730
rect 284354 135702 297836 135716
rect 2137 134526 2142 134554
rect 2170 134526 100044 134554
rect 279972 134526 287686 134554
rect 287714 134526 287719 134554
rect -480 131306 240 131404
rect -480 131292 98686 131306
rect 196 131278 98686 131292
rect 98714 131278 98719 131306
rect 297780 129122 298500 129220
rect 286841 129094 286846 129122
rect 286874 129108 298500 129122
rect 286874 129094 297836 129108
rect 2305 127134 2310 127162
rect 2338 127134 100044 127162
rect 279972 127134 281862 127162
rect 281890 127134 281895 127162
rect 281451 126854 281470 126882
rect 281498 126854 281503 126882
rect -480 124250 240 124348
rect -480 124236 98798 124250
rect 196 124222 98798 124236
rect 98826 124222 98831 124250
rect 297780 122514 298500 122612
rect 281465 122486 281470 122514
rect 281498 122500 298500 122514
rect 281498 122486 297836 122500
rect 98793 119742 98798 119770
rect 98826 119742 100044 119770
rect 279972 119742 282198 119770
rect 282226 119742 282231 119770
rect 281521 119294 281526 119322
rect 281554 119294 282142 119322
rect 282170 119294 282175 119322
rect 196 117292 2198 117306
rect -480 117278 2198 117292
rect 2226 117278 2231 117306
rect -480 117180 240 117278
rect 297780 115962 298500 116004
rect 283481 115934 283486 115962
rect 283514 115934 298500 115962
rect 297780 115892 298500 115934
rect 2193 112350 2198 112378
rect 2226 112350 100044 112378
rect 279972 112350 285166 112378
rect 285194 112350 285199 112378
rect -480 110138 240 110236
rect -480 110124 98966 110138
rect 196 110110 98966 110124
rect 98994 110110 98999 110138
rect 297780 109298 298500 109396
rect 286001 109270 286006 109298
rect 286034 109284 298500 109298
rect 286034 109270 297836 109284
rect 2361 104958 2366 104986
rect 2394 104958 100044 104986
rect 279972 104958 281750 104986
rect 281778 104958 281783 104986
rect 281577 104902 281582 104930
rect 281610 104902 282198 104930
rect 282226 104902 282231 104930
rect -480 103082 240 103180
rect -480 103068 98910 103082
rect 196 103054 98910 103068
rect 98938 103054 98943 103082
rect 297780 102690 298500 102788
rect 282137 102662 282142 102690
rect 282170 102676 298500 102690
rect 282170 102662 297836 102676
rect 142417 99078 142422 99106
rect 142450 99078 143486 99106
rect 143514 99078 143519 99106
rect 155857 99078 155862 99106
rect 155890 99078 156926 99106
rect 156954 99078 156959 99106
rect 157537 99078 157542 99106
rect 157570 99078 159166 99106
rect 159194 99078 159199 99106
rect 170977 99078 170982 99106
rect 171010 99078 172046 99106
rect 172074 99078 172079 99106
rect 172657 99078 172662 99106
rect 172690 99078 173726 99106
rect 173754 99078 173759 99106
rect 176017 99078 176022 99106
rect 176050 99078 176526 99106
rect 176554 99078 176559 99106
rect 179377 99078 179382 99106
rect 179410 99078 179886 99106
rect 179914 99078 179919 99106
rect 195281 99078 195286 99106
rect 195314 99078 196686 99106
rect 196714 99078 196719 99106
rect 198641 99078 198646 99106
rect 198674 99078 202846 99106
rect 202874 99078 202879 99106
rect 216393 99078 216398 99106
rect 216426 99078 217966 99106
rect 217994 99078 217999 99106
rect 228097 99078 228102 99106
rect 228130 99078 233086 99106
rect 233114 99078 233119 99106
rect 233529 99078 233534 99106
rect 233562 99078 234766 99106
rect 234794 99078 234799 99106
rect 240809 99078 240814 99106
rect 240842 99078 244286 99106
rect 244314 99078 244319 99106
rect 245569 99078 245574 99106
rect 245602 99078 247086 99106
rect 247114 99078 247119 99106
rect 247473 99078 247478 99106
rect 247506 99078 248206 99106
rect 248234 99078 248239 99106
rect 251561 99078 251566 99106
rect 251594 99078 253190 99106
rect 253218 99078 253223 99106
rect 256041 99078 256046 99106
rect 256074 99078 256662 99106
rect 256690 99078 256695 99106
rect 257721 99078 257726 99106
rect 257754 99078 258342 99106
rect 258370 99078 258375 99106
rect 261641 99078 261646 99106
rect 261674 99078 262486 99106
rect 262514 99078 262519 99106
rect 264441 99078 264446 99106
rect 264474 99078 265398 99106
rect 265426 99078 265431 99106
rect 265561 99078 265566 99106
rect 265594 99078 266742 99106
rect 266770 99078 266775 99106
rect 154177 99022 154182 99050
rect 154210 99022 156366 99050
rect 156394 99022 156399 99050
rect 169297 99022 169302 99050
rect 169330 99022 173166 99050
rect 173194 99022 173199 99050
rect 239857 99022 239862 99050
rect 239890 99022 243726 99050
rect 243754 99022 243759 99050
rect 246577 99022 246582 99050
rect 246610 99022 247646 99050
rect 247674 99022 247679 99050
rect 252121 99022 252126 99050
rect 252154 99022 254142 99050
rect 254170 99022 254175 99050
rect 263881 99022 263886 99050
rect 263914 99022 265062 99050
rect 265090 99022 265095 99050
rect 139057 98966 139062 98994
rect 139090 98966 141806 98994
rect 141834 98966 141839 98994
rect 174337 98966 174342 98994
rect 174370 98966 177646 98994
rect 177674 98966 177679 98994
rect 253241 98966 253246 98994
rect 253274 98966 255990 98994
rect 256018 98966 256023 98994
rect 104561 98910 104566 98938
rect 104594 98910 150206 98938
rect 150234 98910 150239 98938
rect 105793 98854 105798 98882
rect 105826 98854 165326 98882
rect 165354 98854 165359 98882
rect 177641 98854 177646 98882
rect 177674 98854 183246 98882
rect 183274 98854 183279 98882
rect 96161 98798 96166 98826
rect 96194 98798 158606 98826
rect 158634 98798 158639 98826
rect 165937 98798 165942 98826
rect 165970 98798 182126 98826
rect 182154 98798 182159 98826
rect 184417 98798 184422 98826
rect 184450 98798 187726 98826
rect 187754 98798 187759 98826
rect 207937 98798 207942 98826
rect 207970 98798 216286 98826
rect 216314 98798 216319 98826
rect 228489 98798 228494 98826
rect 228522 98798 237006 98826
rect 237034 98798 237039 98826
rect 262761 98798 262766 98826
rect 262794 98798 270102 98826
rect 270130 98798 270135 98826
rect 58361 98742 58366 98770
rect 58394 98742 131726 98770
rect 131754 98742 131759 98770
rect 159161 98742 159166 98770
rect 159194 98742 195566 98770
rect 195594 98742 195599 98770
rect 199537 98742 199542 98770
rect 199570 98742 214046 98770
rect 214074 98742 214079 98770
rect 214657 98742 214662 98770
rect 214690 98742 219646 98770
rect 219674 98742 219679 98770
rect 222721 98742 222726 98770
rect 222754 98742 233646 98770
rect 233674 98742 233679 98770
rect 255481 98742 255486 98770
rect 255514 98742 259854 98770
rect 259882 98742 259887 98770
rect 267801 98742 267806 98770
rect 267834 98742 275926 98770
rect 275954 98742 275959 98770
rect 5665 98686 5670 98714
rect 5698 98686 105966 98714
rect 105994 98686 105999 98714
rect 135697 98686 135702 98714
rect 135730 98686 141246 98714
rect 141274 98686 141279 98714
rect 145721 98686 145726 98714
rect 145754 98686 186606 98714
rect 186634 98686 186639 98714
rect 187721 98686 187726 98714
rect 187754 98686 188846 98714
rect 188874 98686 188879 98714
rect 191137 98686 191142 98714
rect 191170 98686 212366 98714
rect 212394 98686 212399 98714
rect 216281 98686 216286 98714
rect 216314 98686 229166 98714
rect 229194 98686 229199 98714
rect 234145 98686 234150 98714
rect 234178 98686 240366 98714
rect 240394 98686 240399 98714
rect 256601 98686 256606 98714
rect 256634 98686 261758 98714
rect 261786 98686 261791 98714
rect 266121 98686 266126 98714
rect 266154 98686 277942 98714
rect 277970 98686 277975 98714
rect 253801 98406 253806 98434
rect 253834 98406 257054 98434
rect 257082 98406 257087 98434
rect 194497 98350 194502 98378
rect 194530 98350 198926 98378
rect 198954 98350 198959 98378
rect 243665 98350 243670 98378
rect 243698 98350 245966 98378
rect 245994 98350 245999 98378
rect 251001 98350 251006 98378
rect 251034 98350 252238 98378
rect 252266 98350 252271 98378
rect 124273 98294 124278 98322
rect 124306 98294 128366 98322
rect 128394 98294 128399 98322
rect 137377 98294 137382 98322
rect 137410 98294 140686 98322
rect 140714 98294 140719 98322
rect 186097 98294 186102 98322
rect 186130 98294 187166 98322
rect 187194 98294 187199 98322
rect 221377 98294 221382 98322
rect 221410 98294 223006 98322
rect 223034 98294 223039 98322
rect 244617 98294 244622 98322
rect 244650 98294 246526 98322
rect 246554 98294 246559 98322
rect 250441 98294 250446 98322
rect 250474 98294 251286 98322
rect 251314 98294 251319 98322
rect 86585 97902 86590 97930
rect 86618 97902 153566 97930
rect 153594 97902 153599 97930
rect 265393 97902 265398 97930
rect 265426 97902 275086 97930
rect 275114 97902 275119 97930
rect 11377 97846 11382 97874
rect 11410 97846 109326 97874
rect 109354 97846 109359 97874
rect 147513 97846 147518 97874
rect 147546 97846 189406 97874
rect 189434 97846 189439 97874
rect 226529 97846 226534 97874
rect 226562 97846 235886 97874
rect 235914 97846 235919 97874
rect 271161 97846 271166 97874
rect 271194 97846 286510 97874
rect 286538 97846 286543 97874
rect 68497 97062 68502 97090
rect 68530 97062 142758 97090
rect 142786 97062 142791 97090
rect 15185 97006 15190 97034
rect 15218 97006 111566 97034
rect 111594 97006 111599 97034
rect 117049 97006 117054 97034
rect 117082 97006 171318 97034
rect 171346 97006 171351 97034
rect 224625 97006 224630 97034
rect 224658 97006 233534 97034
rect 233562 97006 233567 97034
rect 269481 97006 269486 97034
rect 269514 97006 283654 97034
rect 283682 97006 283687 97034
rect 98009 96222 98014 96250
rect 98042 96222 160286 96250
rect 160314 96222 160319 96250
rect 43745 96166 43750 96194
rect 43778 96166 124278 96194
rect 124306 96166 124311 96194
rect 270041 96166 270046 96194
rect 270074 96166 284606 96194
rect 284634 96166 284639 96194
rect 196 96124 3766 96138
rect -480 96110 3766 96124
rect 3794 96110 3799 96138
rect -480 96012 240 96110
rect 297780 96082 298500 96180
rect 282641 96054 282646 96082
rect 282674 96068 298500 96082
rect 282674 96054 297836 96068
rect 103721 93702 103726 93730
rect 103754 93702 163646 93730
rect 163674 93702 163679 93730
rect 46601 93646 46606 93674
rect 46634 93646 130046 93674
rect 130074 93646 130079 93674
rect 266737 93646 266742 93674
rect 266770 93646 276990 93674
rect 277018 93646 277023 93674
rect 91345 92862 91350 92890
rect 91378 92862 154182 92890
rect 154210 92862 154215 92890
rect 52313 92806 52318 92834
rect 52346 92806 133406 92834
rect 133434 92806 133439 92834
rect 94201 91182 94206 91210
rect 94234 91182 157654 91210
rect 157682 91182 157687 91210
rect 55169 91126 55174 91154
rect 55202 91126 135086 91154
rect 135114 91126 135119 91154
rect 66593 90286 66598 90314
rect 66626 90286 139062 90314
rect 139090 90286 139095 90314
rect 292721 89558 292726 89586
rect 292754 89572 297836 89586
rect 292754 89558 298500 89572
rect 69449 89446 69454 89474
rect 69482 89446 142422 89474
rect 142450 89446 142455 89474
rect 297780 89460 298500 89558
rect -480 88970 240 89068
rect -480 88956 99022 88970
rect 196 88942 99022 88956
rect 99050 88942 99055 88970
rect 89441 88606 89446 88634
rect 89474 88606 155246 88634
rect 155274 88606 155279 88634
rect 72305 87766 72310 87794
rect 72338 87766 145166 87794
rect 145194 87766 145199 87794
rect 75161 86982 75166 87010
rect 75194 86982 146846 87010
rect 146874 86982 146879 87010
rect 24705 86926 24710 86954
rect 24738 86926 117166 86954
rect 117194 86926 117199 86954
rect 78017 85246 78022 85274
rect 78050 85246 148526 85274
rect 148554 85246 148559 85274
rect 83729 84462 83734 84490
rect 83762 84462 151886 84490
rect 151914 84462 151919 84490
rect 17089 84406 17094 84434
rect 17122 84406 112686 84434
rect 112714 84406 112719 84434
rect 297780 82866 298500 82964
rect 282193 82838 282198 82866
rect 282226 82852 298500 82866
rect 282226 82838 297836 82852
rect -480 81914 240 82012
rect -480 81900 98630 81914
rect 196 81886 98630 81900
rect 98658 81886 98663 81914
rect 100865 81886 100870 81914
rect 100898 81886 161966 81914
rect 161994 81886 161999 81914
rect 92297 81102 92302 81130
rect 92330 81102 155862 81130
rect 155890 81102 155895 81130
rect 21401 81046 21406 81074
rect 21434 81046 114366 81074
rect 114394 81046 114399 81074
rect 22801 80206 22806 80234
rect 22834 80206 116046 80234
rect 116074 80206 116079 80234
rect 26609 79366 26614 79394
rect 26642 79366 118286 79394
rect 118314 79366 118319 79394
rect 29465 78526 29470 78554
rect 29498 78526 119966 78554
rect 119994 78526 119999 78554
rect 32321 77686 32326 77714
rect 32354 77686 121646 77714
rect 121674 77686 121679 77714
rect 297780 76258 298500 76356
rect 281913 76230 281918 76258
rect 281946 76244 298500 76258
rect 281946 76230 297836 76244
rect 35177 76006 35182 76034
rect 35210 76006 123326 76034
rect 123354 76006 123359 76034
rect 177977 76006 177982 76034
rect 178010 76006 207326 76034
rect 207354 76006 207359 76034
rect 38033 75166 38038 75194
rect 38066 75166 125006 75194
rect 125034 75166 125039 75194
rect 196 74956 2254 74970
rect -480 74942 2254 74956
rect 2282 74942 2287 74970
rect -480 74844 240 74942
rect 64689 72646 64694 72674
rect 64722 72646 137382 72674
rect 137410 72646 137415 72674
rect 73257 71806 73262 71834
rect 73290 71806 145670 71834
rect 145698 71806 145703 71834
rect 76113 70966 76118 70994
rect 76146 70966 147406 70994
rect 147434 70966 147439 70994
rect 62785 70126 62790 70154
rect 62818 70126 139566 70154
rect 139594 70126 139599 70154
rect 297780 69650 298500 69748
rect 289361 69622 289366 69650
rect 289394 69636 298500 69650
rect 289394 69622 297836 69636
rect 101817 69286 101822 69314
rect 101850 69286 162526 69314
rect 162554 69286 162559 69314
rect 162745 69286 162750 69314
rect 162778 69286 198366 69314
rect 198394 69286 198399 69314
rect -480 67802 240 67900
rect -480 67788 99078 67802
rect 196 67774 99078 67788
rect 99106 67774 99111 67802
rect 39937 66766 39942 66794
rect 39970 66766 126126 66794
rect 126154 66766 126159 66794
rect 154177 65982 154182 66010
rect 154210 65982 193326 66010
rect 193354 65982 193359 66010
rect 87537 65926 87542 65954
rect 87570 65926 154126 65954
rect 154154 65926 154159 65954
rect 42849 64246 42854 64274
rect 42882 64246 127806 64274
rect 127834 64246 127839 64274
rect 143705 64246 143710 64274
rect 143738 64246 186102 64274
rect 186130 64246 186135 64274
rect 297780 63042 298500 63140
rect 281969 63014 281974 63042
rect 282002 63028 298500 63042
rect 282002 63014 297836 63028
rect 14289 61726 14294 61754
rect 14322 61726 111006 61754
rect 111034 61726 111039 61754
rect -480 60746 240 60844
rect -480 60732 98686 60746
rect 196 60718 98686 60732
rect 98714 60718 98719 60746
rect 88489 60046 88494 60074
rect 88522 60046 154686 60074
rect 154714 60046 154719 60074
rect 51361 58366 51366 58394
rect 51394 58366 132846 58394
rect 132874 58366 132879 58394
rect 67545 57526 67550 57554
rect 67578 57526 142366 57554
rect 142394 57526 142399 57554
rect 56121 56686 56126 56714
rect 56154 56686 135646 56714
rect 135674 56686 135679 56714
rect 297780 56434 298500 56532
rect 282025 56406 282030 56434
rect 282058 56420 298500 56434
rect 282058 56406 297836 56420
rect 47553 55006 47558 55034
rect 47586 55006 130606 55034
rect 130634 55006 130639 55034
rect 18993 54166 18998 54194
rect 19026 54166 113806 54194
rect 113834 54166 113839 54194
rect -480 53746 240 53788
rect -480 53718 2086 53746
rect 2114 53718 2119 53746
rect -480 53676 240 53718
rect 82777 53326 82782 53354
rect 82810 53326 151326 53354
rect 151354 53326 151359 53354
rect 23753 52486 23758 52514
rect 23786 52486 116606 52514
rect 116634 52486 116639 52514
rect 93249 51646 93254 51674
rect 93282 51646 157486 51674
rect 157514 51646 157519 51674
rect 258281 51646 258286 51674
rect 258314 51646 264614 51674
rect 264642 51646 264647 51674
rect 265057 51646 265062 51674
rect 265090 51646 274134 51674
rect 274162 51646 274167 51674
rect 297780 49826 298500 49924
rect 282081 49798 282086 49826
rect 282114 49812 298500 49826
rect 282114 49798 297836 49812
rect 37081 48286 37086 48314
rect 37114 48286 124446 48314
rect 124474 48286 124479 48314
rect -480 46634 240 46732
rect -480 46620 98742 46634
rect 196 46606 98742 46620
rect 98770 46606 98775 46634
rect 61833 44926 61838 44954
rect 61866 44926 139006 44954
rect 139034 44926 139039 44954
rect 85689 44086 85694 44114
rect 85722 44086 153006 44114
rect 153034 44086 153039 44114
rect 268921 44086 268926 44114
rect 268954 44086 282702 44114
rect 282730 44086 282735 44114
rect 48505 43246 48510 43274
rect 48538 43246 131166 43274
rect 131194 43246 131199 43274
rect 297780 43218 298500 43316
rect 282137 43190 282142 43218
rect 282170 43204 298500 43218
rect 282170 43190 297836 43204
rect 31369 42406 31374 42434
rect 31402 42406 121086 42434
rect 121114 42406 121119 42434
rect 200825 42406 200830 42434
rect 200858 42406 220766 42434
rect 220794 42406 220799 42434
rect 102769 39886 102774 39914
rect 102802 39886 163086 39914
rect 163114 39886 163119 39914
rect -480 39578 240 39676
rect -480 39564 98854 39578
rect 196 39550 98854 39564
rect 98882 39550 98887 39578
rect 99969 39046 99974 39074
rect 100002 39046 161406 39074
rect 161434 39046 161439 39074
rect 77065 37366 77070 37394
rect 77098 37366 147966 37394
rect 147994 37366 147999 37394
rect 297780 36610 298500 36708
rect 281801 36582 281806 36610
rect 281834 36596 298500 36610
rect 281834 36582 297836 36596
rect 90393 36526 90398 36554
rect 90426 36526 155806 36554
rect 155834 36526 155839 36554
rect 104673 35686 104678 35714
rect 104706 35686 164206 35714
rect 164234 35686 164239 35714
rect 53265 34846 53270 34874
rect 53298 34846 133966 34874
rect 133994 34846 133999 34874
rect 128529 34062 128534 34090
rect 128562 34062 178206 34090
rect 178234 34062 178239 34090
rect 44697 34006 44702 34034
rect 44730 34006 128926 34034
rect 128954 34006 128959 34034
rect 30417 33166 30422 33194
rect 30450 33166 120526 33194
rect 120554 33166 120559 33194
rect 134185 33166 134190 33194
rect 134218 33166 181566 33194
rect 181594 33166 181599 33194
rect 196 32620 2142 32634
rect -480 32606 2142 32620
rect 2170 32606 2175 32634
rect -480 32508 240 32606
rect 137041 30702 137046 30730
rect 137074 30702 177646 30730
rect 177674 30702 177679 30730
rect 58977 30646 58982 30674
rect 59010 30646 137326 30674
rect 137354 30646 137359 30674
rect 297780 30002 298500 30100
rect 287681 29974 287686 30002
rect 287714 29988 298500 30002
rect 287714 29974 297836 29988
rect 108481 29806 108486 29834
rect 108514 29806 166446 29834
rect 166474 29806 166479 29834
rect 183521 29806 183526 29834
rect 183554 29806 210126 29834
rect 210154 29806 210159 29834
rect 28569 28126 28574 28154
rect 28602 28126 119406 28154
rect 119434 28126 119439 28154
rect 130377 28126 130382 28154
rect 130410 28126 179326 28154
rect 179354 28126 179359 28154
rect 182849 28126 182854 28154
rect 182882 28126 208446 28154
rect 208474 28126 208479 28154
rect 172713 27342 172718 27370
rect 172746 27342 203406 27370
rect 203434 27342 203439 27370
rect 6617 27286 6622 27314
rect 6650 27286 106526 27314
rect 106554 27286 106559 27314
rect 121809 27286 121814 27314
rect 121842 27286 174286 27314
rect 174314 27286 174319 27314
rect 267241 27286 267246 27314
rect 267274 27286 279846 27314
rect 279874 27286 279879 27314
rect 168457 26502 168462 26530
rect 168490 26502 201726 26530
rect 201754 26502 201759 26530
rect 27561 26446 27566 26474
rect 27594 26446 118846 26474
rect 118874 26446 118879 26474
rect 118953 26446 118958 26474
rect 118986 26446 172606 26474
rect 172634 26446 172639 26474
rect 157089 25662 157094 25690
rect 157122 25662 195006 25690
rect 195034 25662 195039 25690
rect 116097 25606 116102 25634
rect 116130 25606 170926 25634
rect 170954 25606 170959 25634
rect 197017 25606 197022 25634
rect 197050 25606 218526 25634
rect 218554 25606 218559 25634
rect 196 25564 2310 25578
rect -480 25550 2310 25564
rect 2338 25550 2343 25578
rect -480 25452 240 25550
rect 156081 24822 156086 24850
rect 156114 24822 194446 24850
rect 194474 24822 194479 24850
rect 111337 24766 111342 24794
rect 111370 24766 168126 24794
rect 168154 24766 168159 24794
rect 195337 24766 195342 24794
rect 195370 24766 216846 24794
rect 216874 24766 216879 24794
rect 150369 23982 150374 24010
rect 150402 23982 191086 24010
rect 191114 23982 191119 24010
rect 114249 23926 114254 23954
rect 114282 23926 169806 23954
rect 169834 23926 169839 23954
rect 192817 23926 192822 23954
rect 192850 23926 215166 23954
rect 215194 23926 215199 23954
rect 297780 23394 298500 23492
rect 281857 23366 281862 23394
rect 281890 23380 298500 23394
rect 281890 23366 297836 23380
rect 138945 22302 138950 22330
rect 138978 22302 184366 22330
rect 184394 22302 184399 22330
rect 96105 22246 96110 22274
rect 96138 22246 157542 22274
rect 157570 22246 157575 22274
rect 185649 22246 185654 22274
rect 185682 22246 211806 22274
rect 211834 22246 211839 22274
rect 132337 21462 132342 21490
rect 132370 21462 180446 21490
rect 180474 21462 180479 21490
rect 105625 21406 105630 21434
rect 105658 21406 164766 21434
rect 164794 21406 164799 21434
rect 174169 21406 174174 21434
rect 174202 21406 205086 21434
rect 205114 21406 205119 21434
rect 207041 21406 207046 21434
rect 207074 21406 223566 21434
rect 223594 21406 223599 21434
rect 262201 21406 262206 21434
rect 262234 21406 271334 21434
rect 271362 21406 271367 21434
rect 129425 18942 129430 18970
rect 129458 18942 178766 18970
rect 178794 18942 178799 18970
rect 81825 18886 81830 18914
rect 81858 18886 150766 18914
rect 150794 18886 150799 18914
rect 151321 18886 151326 18914
rect 151354 18886 191646 18914
rect 191674 18886 191679 18914
rect 196065 18886 196070 18914
rect 196098 18886 216398 18914
rect 216426 18886 216431 18914
rect -480 18410 240 18508
rect -480 18396 98798 18410
rect 196 18382 98798 18396
rect 98826 18382 98831 18410
rect 126569 18102 126574 18130
rect 126602 18102 177086 18130
rect 177114 18102 177119 18130
rect 98961 18046 98966 18074
rect 98994 18046 160846 18074
rect 160874 18046 160879 18074
rect 178929 18046 178934 18074
rect 178962 18046 207886 18074
rect 207914 18046 207919 18074
rect 119905 17262 119910 17290
rect 119938 17262 169302 17290
rect 169330 17262 169335 17290
rect 170417 17262 170422 17290
rect 170450 17262 198646 17290
rect 198674 17262 198679 17290
rect 123713 17206 123718 17234
rect 123746 17206 175406 17234
rect 175434 17206 175439 17234
rect 177025 17206 177030 17234
rect 177058 17206 206766 17234
rect 206794 17206 206799 17234
rect 297780 16842 298500 16884
rect 282193 16814 282198 16842
rect 282226 16814 298500 16842
rect 297780 16772 298500 16814
rect 131329 16422 131334 16450
rect 131362 16422 179382 16450
rect 179410 16422 179415 16450
rect 113297 16366 113302 16394
rect 113330 16366 169246 16394
rect 169274 16366 169279 16394
rect 169409 16366 169414 16394
rect 169442 16366 202286 16394
rect 202314 16366 202319 16394
rect 203737 16366 203742 16394
rect 203770 16366 221886 16394
rect 221914 16366 221919 16394
rect 120857 15582 120862 15610
rect 120890 15582 172662 15610
rect 172690 15582 172695 15610
rect 180833 15582 180838 15610
rect 180866 15582 209006 15610
rect 209034 15582 209039 15610
rect 34225 15526 34230 15554
rect 34258 15526 122766 15554
rect 122794 15526 122799 15554
rect 133233 15526 133238 15554
rect 133266 15526 181006 15554
rect 181034 15526 181039 15554
rect 148465 14742 148470 14770
rect 148498 14742 189966 14770
rect 189994 14742 189999 14770
rect 190241 14742 190246 14770
rect 190274 14742 213486 14770
rect 213514 14742 213519 14770
rect 20897 14686 20902 14714
rect 20930 14686 114926 14714
rect 114954 14686 114959 14714
rect 115145 14686 115150 14714
rect 115178 14686 170366 14714
rect 170394 14686 170399 14714
rect 172265 14686 172270 14714
rect 172298 14686 203966 14714
rect 203994 14686 203999 14714
rect 166553 13118 166558 13146
rect 166586 13118 200606 13146
rect 200634 13118 200639 13146
rect 109433 13062 109438 13090
rect 109466 13062 167006 13090
rect 167034 13062 167039 13090
rect 50409 13006 50414 13034
rect 50442 13006 132286 13034
rect 132314 13006 132319 13034
rect 145609 13006 145614 13034
rect 145642 13006 188286 13034
rect 188314 13006 188319 13034
rect 201777 13006 201782 13034
rect 201810 13006 221326 13034
rect 221354 13006 221359 13034
rect 165601 12278 165606 12306
rect 165634 12278 200046 12306
rect 200074 12278 200079 12306
rect 80873 12222 80878 12250
rect 80906 12222 104566 12250
rect 104594 12222 104599 12250
rect 118001 12222 118006 12250
rect 118034 12222 170982 12250
rect 171010 12222 171015 12250
rect 213201 12222 213206 12250
rect 213234 12222 228046 12250
rect 228074 12222 228079 12250
rect 65641 12166 65646 12194
rect 65674 12166 135702 12194
rect 135730 12166 135735 12194
rect 160841 12166 160846 12194
rect 160874 12166 197246 12194
rect 197274 12166 197279 12194
rect 198921 12166 198926 12194
rect 198954 12166 214662 12194
rect 214690 12166 214695 12194
rect 196 11452 2198 11466
rect -480 11438 2198 11452
rect 2226 11438 2231 11466
rect -480 11340 240 11438
rect 159889 10542 159894 10570
rect 159922 10542 195286 10570
rect 195314 10542 195319 10570
rect 124665 10486 124670 10514
rect 124698 10486 175966 10514
rect 175994 10486 175999 10514
rect 199929 10486 199934 10514
rect 199962 10486 220206 10514
rect 220234 10486 220239 10514
rect 297780 10178 298500 10276
rect 285161 10150 285166 10178
rect 285194 10164 298500 10178
rect 285194 10150 297836 10164
rect 161793 9758 161798 9786
rect 161826 9758 197806 9786
rect 197834 9758 197839 9786
rect 78969 9702 78974 9730
rect 79002 9702 149086 9730
rect 149114 9702 149119 9730
rect 149417 9702 149422 9730
rect 149450 9702 190526 9730
rect 190554 9702 190559 9730
rect 210345 9702 210350 9730
rect 210378 9702 226366 9730
rect 226394 9702 226399 9730
rect 7569 9646 7574 9674
rect 7602 9646 107086 9674
rect 107114 9646 107119 9674
rect 107529 9646 107534 9674
rect 107562 9646 165886 9674
rect 165914 9646 165919 9674
rect 187497 9646 187502 9674
rect 187530 9646 212926 9674
rect 212954 9646 212959 9674
rect 144657 8974 144662 9002
rect 144690 8974 184422 9002
rect 184450 8974 184455 9002
rect 79921 8918 79926 8946
rect 79954 8918 149646 8946
rect 149674 8918 149679 8946
rect 74209 8862 74214 8890
rect 74242 8862 146286 8890
rect 146314 8862 146319 8890
rect 184641 8862 184646 8890
rect 184674 8862 211246 8890
rect 211274 8862 211279 8890
rect 71409 8806 71414 8834
rect 71442 8806 144606 8834
rect 144634 8806 144639 8834
rect 155129 8806 155134 8834
rect 155162 8806 193886 8834
rect 193914 8806 193919 8834
rect 203681 8806 203686 8834
rect 203714 8806 222446 8834
rect 222474 8806 222479 8834
rect 59929 8078 59934 8106
rect 59962 8078 137886 8106
rect 137914 8078 137919 8106
rect 183689 8078 183694 8106
rect 183722 8078 210686 8106
rect 210714 8078 210719 8106
rect 57129 8022 57134 8050
rect 57162 8022 136206 8050
rect 136234 8022 136239 8050
rect 153225 8022 153230 8050
rect 153258 8022 192766 8050
rect 192794 8022 192799 8050
rect 193209 8022 193214 8050
rect 193242 8022 207942 8050
rect 207970 8022 207975 8050
rect 54217 7966 54222 7994
rect 54250 7966 134526 7994
rect 134554 7966 134559 7994
rect 137993 7966 137998 7994
rect 138026 7966 183806 7994
rect 183834 7966 183839 7994
rect 207489 7966 207494 7994
rect 207522 7966 224686 7994
rect 224714 7966 224719 7994
rect 265001 7966 265006 7994
rect 265034 7966 276038 7994
rect 276066 7966 276071 7994
rect 84681 7238 84686 7266
rect 84714 7238 152446 7266
rect 152474 7238 152479 7266
rect 181785 7238 181790 7266
rect 181818 7238 209566 7266
rect 209594 7238 209599 7266
rect 45649 7182 45654 7210
rect 45682 7182 129486 7210
rect 129514 7182 129519 7210
rect 152273 7182 152278 7210
rect 152306 7182 192206 7210
rect 192234 7182 192239 7210
rect 41841 7126 41846 7154
rect 41874 7126 127246 7154
rect 127274 7126 127279 7154
rect 136089 7126 136094 7154
rect 136122 7126 182686 7154
rect 182714 7126 182719 7154
rect 197969 7126 197974 7154
rect 198002 7126 219086 7154
rect 219114 7126 219119 7154
rect 220817 7126 220822 7154
rect 220850 7126 232526 7154
rect 232554 7126 232559 7154
rect 259961 7126 259966 7154
rect 259994 7126 267470 7154
rect 267498 7126 267503 7154
rect 271721 7126 271726 7154
rect 271754 7126 287462 7154
rect 287490 7126 287495 7154
rect 70401 6398 70406 6426
rect 70434 6398 144046 6426
rect 144074 6398 144079 6426
rect 158937 6398 158942 6426
rect 158970 6398 196126 6426
rect 196154 6398 196159 6426
rect 38985 6342 38990 6370
rect 39018 6342 125566 6370
rect 125594 6342 125599 6370
rect 146561 6342 146566 6370
rect 146594 6342 187726 6370
rect 187754 6342 187759 6370
rect 190353 6342 190358 6370
rect 190386 6342 214606 6370
rect 214634 6342 214639 6370
rect 218913 6342 218918 6370
rect 218946 6342 231406 6370
rect 231434 6342 231439 6370
rect 36129 6286 36134 6314
rect 36162 6286 123886 6314
rect 123914 6286 123919 6314
rect 127521 6286 127526 6314
rect 127554 6286 174342 6314
rect 174370 6286 174375 6314
rect 175121 6286 175126 6314
rect 175154 6286 205646 6314
rect 205674 6286 205679 6314
rect 212249 6286 212254 6314
rect 212282 6286 227486 6314
rect 227514 6286 227519 6314
rect 232241 6286 232246 6314
rect 232274 6286 239246 6314
rect 239274 6286 239279 6314
rect 259401 6286 259406 6314
rect 259434 6286 266518 6314
rect 266546 6286 266551 6314
rect 268361 6286 268366 6314
rect 268394 6286 281750 6314
rect 281778 6286 281783 6314
rect 33385 5446 33390 5474
rect 33418 5446 122206 5474
rect 122234 5446 122239 5474
rect 140009 5446 140014 5474
rect 140042 5446 184926 5474
rect 184954 5446 184959 5474
rect 110497 4718 110502 4746
rect 110530 4718 167566 4746
rect 167594 4718 167599 4746
rect 16249 4662 16254 4690
rect 16282 4662 112126 4690
rect 112154 4662 112159 4690
rect 164761 4662 164766 4690
rect 164794 4662 199486 4690
rect 199514 4662 199519 4690
rect 13393 4606 13398 4634
rect 13426 4606 110446 4634
rect 110474 4606 110479 4634
rect 125729 4606 125734 4634
rect 125762 4606 176022 4634
rect 176050 4606 176055 4634
rect 216169 4606 216174 4634
rect 216202 4606 229726 4634
rect 229754 4606 229759 4634
rect 196 4396 2366 4410
rect -480 4382 2366 4396
rect 2394 4382 2399 4410
rect -480 4284 240 4382
rect 41001 3878 41006 3906
rect 41034 3878 126686 3906
rect 126714 3878 126719 3906
rect 135193 3878 135198 3906
rect 135226 3878 165942 3906
rect 165970 3878 165975 3906
rect 167617 3878 167622 3906
rect 167650 3878 201166 3906
rect 201194 3878 201199 3906
rect 258337 3878 258342 3906
rect 258370 3878 263662 3906
rect 263690 3878 263695 3906
rect 12441 3822 12446 3850
rect 12474 3822 109886 3850
rect 109914 3822 109919 3850
rect 122873 3822 122878 3850
rect 122906 3822 174846 3850
rect 174874 3822 174879 3850
rect 176185 3822 176190 3850
rect 176218 3822 206206 3850
rect 206234 3822 206239 3850
rect 209505 3822 209510 3850
rect 209538 3822 225806 3850
rect 225834 3822 225839 3850
rect 262481 3822 262486 3850
rect 262514 3822 270326 3850
rect 270354 3822 270359 3850
rect 8633 3766 8638 3794
rect 8666 3766 107646 3794
rect 107674 3766 107679 3794
rect 112401 3766 112406 3794
rect 112434 3766 168686 3794
rect 168714 3766 168719 3794
rect 173329 3766 173334 3794
rect 173362 3766 204526 3794
rect 204554 3766 204559 3794
rect 204745 3766 204750 3794
rect 204778 3766 221382 3794
rect 221410 3766 221415 3794
rect 223785 3766 223790 3794
rect 223818 3766 234206 3794
rect 234234 3766 234239 3794
rect 263321 3766 263326 3794
rect 263354 3766 273182 3794
rect 273210 3766 273215 3794
rect 297780 3570 298500 3668
rect 281745 3542 281750 3570
rect 281778 3556 298500 3570
rect 281778 3542 297836 3556
rect 189513 3094 189518 3122
rect 189546 3094 199542 3122
rect 199570 3094 199575 3122
rect 63793 3038 63798 3066
rect 63826 3038 140126 3066
rect 140154 3038 140159 3066
rect 141913 3038 141918 3066
rect 141946 3038 151214 3066
rect 163753 3038 163758 3066
rect 163786 3038 194502 3066
rect 194530 3038 194535 3066
rect 206593 3038 206598 3066
rect 206626 3038 224126 3066
rect 224154 3038 224159 3066
rect 151186 3010 151214 3038
rect 49513 2982 49518 3010
rect 49546 2982 58366 3010
rect 58394 2982 58399 3010
rect 60993 2982 60998 3010
rect 61026 2982 138446 3010
rect 138474 2982 138479 3010
rect 142865 2982 142870 3010
rect 142898 2982 145726 3010
rect 145754 2982 145759 3010
rect 151186 2982 186046 3010
rect 186074 2982 186079 3010
rect 195225 2982 195230 3010
rect 195258 2982 212954 3010
rect 221881 2982 221886 3010
rect 221914 2982 228102 3010
rect 228130 2982 228135 3010
rect 229497 2982 229502 3010
rect 229530 2982 237566 3010
rect 237594 2982 237599 3010
rect 261081 2982 261086 3010
rect 261114 2982 269374 3010
rect 269402 2982 269407 3010
rect 275921 2982 275926 3010
rect 275954 2982 280798 3010
rect 280826 2982 280831 3010
rect 58137 2926 58142 2954
rect 58170 2926 136766 2954
rect 136794 2926 136799 2954
rect 140961 2926 140966 2954
rect 140994 2926 185486 2954
rect 185514 2926 185519 2954
rect 192313 2926 192318 2954
rect 192346 2926 204134 2954
rect 204106 2842 204134 2926
rect 212926 2898 212954 2982
rect 215217 2926 215222 2954
rect 215250 2926 216286 2954
rect 216314 2926 216319 2954
rect 218073 2926 218078 2954
rect 218106 2926 230846 2954
rect 230874 2926 230879 2954
rect 235153 2926 235158 2954
rect 235186 2926 240926 2954
rect 240954 2926 240959 2954
rect 256657 2926 256662 2954
rect 256690 2926 260806 2954
rect 260834 2926 260839 2954
rect 266681 2926 266686 2954
rect 266714 2926 278894 2954
rect 278922 2926 278927 2954
rect 212926 2870 217406 2898
rect 217434 2870 217439 2898
rect 204106 2814 215726 2842
rect 215754 2814 215759 2842
rect 95265 2534 95270 2562
rect 95298 2534 96166 2562
rect 96194 2534 96199 2562
rect 105793 2534 105798 2562
rect 105826 2534 106582 2562
rect 106610 2534 106615 2562
rect 158097 2534 158102 2562
rect 158130 2534 159166 2562
rect 159194 2534 159199 2562
rect 186657 2534 186662 2562
rect 186690 2534 191142 2562
rect 191170 2534 191175 2562
rect 270097 2534 270102 2562
rect 270130 2534 272230 2562
rect 272258 2534 272263 2562
rect 191417 2478 191422 2506
rect 191450 2478 192822 2506
rect 192850 2478 192855 2506
rect 242825 2478 242830 2506
rect 242858 2478 245406 2506
rect 245434 2478 245439 2506
rect 254361 2478 254366 2506
rect 254394 2478 257950 2506
rect 257978 2478 257983 2506
rect 238065 2366 238070 2394
rect 238098 2366 242606 2394
rect 242634 2366 242639 2394
rect 25769 2310 25774 2338
rect 25802 2310 117726 2338
rect 117754 2310 117759 2338
rect 219977 2310 219982 2338
rect 220010 2310 231966 2338
rect 231994 2310 231999 2338
rect 233305 2310 233310 2338
rect 233338 2310 239806 2338
rect 239834 2310 239839 2338
rect 270601 2310 270606 2338
rect 270634 2310 285614 2338
rect 285642 2310 285647 2338
rect 21961 2254 21966 2282
rect 21994 2254 115486 2282
rect 115514 2254 115519 2282
rect 217121 2254 217126 2282
rect 217154 2254 230286 2282
rect 230314 2254 230319 2282
rect 231401 2254 231406 2282
rect 231434 2254 238686 2282
rect 238714 2254 238719 2282
rect 272281 2254 272286 2282
rect 272314 2254 288414 2282
rect 288442 2254 288447 2282
rect 18153 2198 18158 2226
rect 18186 2198 113246 2226
rect 113274 2198 113279 2226
rect 214265 2198 214270 2226
rect 214298 2198 228606 2226
rect 228634 2198 228639 2226
rect 230449 2198 230454 2226
rect 230482 2198 238126 2226
rect 238154 2198 238159 2226
rect 239017 2198 239022 2226
rect 239050 2198 243166 2226
rect 243194 2198 243199 2226
rect 272841 2198 272846 2226
rect 272874 2198 290318 2226
rect 290346 2198 290351 2226
rect 10537 2142 10542 2170
rect 10570 2142 108766 2170
rect 108794 2142 108799 2170
rect 180586 2142 182798 2170
rect 182826 2142 182831 2170
rect 211409 2142 211414 2170
rect 211442 2142 226926 2170
rect 226954 2142 226959 2170
rect 227593 2142 227598 2170
rect 227626 2142 236446 2170
rect 236474 2142 236479 2170
rect 237113 2142 237118 2170
rect 237146 2142 242046 2170
rect 242074 2142 242079 2170
rect 252681 2142 252686 2170
rect 252714 2142 255094 2170
rect 255122 2142 255127 2170
rect 258841 2142 258846 2170
rect 258874 2142 265566 2170
rect 265594 2142 265599 2170
rect 273401 2142 273406 2170
rect 273434 2142 291270 2170
rect 291298 2142 291303 2170
rect 180586 2114 180614 2142
rect 9585 2086 9590 2114
rect 9618 2086 108206 2114
rect 108234 2086 108239 2114
rect 171425 2086 171430 2114
rect 171458 2086 172718 2114
rect 172746 2086 172751 2114
rect 179993 2086 179998 2114
rect 180026 2086 180614 2114
rect 182849 2086 182854 2114
rect 182882 2086 183526 2114
rect 183554 2086 183559 2114
rect 188561 2086 188566 2114
rect 188594 2086 190246 2114
rect 190274 2086 190279 2114
rect 194273 2086 194278 2114
rect 194306 2086 195342 2114
rect 195370 2086 195375 2114
rect 202841 2086 202846 2114
rect 202874 2086 203742 2114
rect 203770 2086 203775 2114
rect 205697 2086 205702 2114
rect 205730 2086 207046 2114
rect 207074 2086 207079 2114
rect 208553 2086 208558 2114
rect 208586 2086 225246 2114
rect 225274 2086 225279 2114
rect 225689 2086 225694 2114
rect 225722 2086 235326 2114
rect 235354 2086 235359 2114
rect 236161 2086 236166 2114
rect 236194 2086 241486 2114
rect 241514 2086 241519 2114
rect 241873 2086 241878 2114
rect 241906 2086 244846 2114
rect 244874 2086 244879 2114
rect 249881 2086 249886 2114
rect 249914 2086 250334 2114
rect 250362 2086 250367 2114
rect 254921 2086 254926 2114
rect 254954 2086 258902 2114
rect 258930 2086 258935 2114
rect 260521 2086 260526 2114
rect 260554 2086 268422 2114
rect 268450 2086 268455 2114
rect 273961 2086 273966 2114
rect 273994 2086 292222 2114
rect 292250 2086 292255 2114
rect 20057 2030 20062 2058
rect 20090 2030 21406 2058
rect 21434 2030 21439 2058
rect 257161 2030 257166 2058
rect 257194 2030 262710 2058
rect 262738 2030 262743 2058
rect 97169 1246 97174 1274
rect 97202 1246 159726 1274
rect 159754 1246 159759 1274
<< via3 >>
rect 98686 274974 98714 275002
rect 281414 274974 281442 275002
rect 2086 267582 2114 267610
rect 281806 267582 281834 267610
rect 98742 260190 98770 260218
rect 281862 260190 281890 260218
rect 98854 252798 98882 252826
rect 284326 252798 284354 252826
rect 2142 245406 2170 245434
rect 286846 245406 286874 245434
rect 281470 238014 281498 238042
rect 98798 230622 98826 230650
rect 283486 230622 283514 230650
rect 2198 223230 2226 223258
rect 286006 223230 286034 223258
rect 98966 215838 98994 215866
rect 281526 215838 281554 215866
rect 98910 208446 98938 208474
rect 282646 208446 282674 208474
rect 3766 201054 3794 201082
rect 292726 201054 292754 201082
rect 99022 193662 99050 193690
rect 281582 193662 281610 193690
rect 98630 186270 98658 186298
rect 281918 186270 281946 186298
rect 2254 178878 2282 178906
rect 289366 178878 289394 178906
rect 99078 171486 99106 171514
rect 281974 171486 282002 171514
rect 98686 166558 98714 166586
rect 98686 164094 98714 164122
rect 282030 164094 282058 164122
rect 2086 159558 2114 159586
rect 2086 156702 2114 156730
rect 282086 156702 282114 156730
rect 281414 156310 281442 156338
rect 98742 152446 98770 152474
rect 98742 149310 98770 149338
rect 282142 149310 282170 149338
rect 281806 148918 281834 148946
rect 98854 145390 98882 145418
rect 281862 142310 281890 142338
rect 98854 141918 98882 141946
rect 281806 141918 281834 141946
rect 2142 138446 2170 138474
rect 284326 135702 284354 135730
rect 2142 134526 2170 134554
rect 287686 134526 287714 134554
rect 286846 129094 286874 129122
rect 2310 127134 2338 127162
rect 281862 127134 281890 127162
rect 281470 126854 281498 126882
rect 98798 124222 98826 124250
rect 98798 119742 98826 119770
rect 282198 119742 282226 119770
rect 281526 119294 281554 119322
rect 2198 117278 2226 117306
rect 283486 115934 283514 115962
rect 2198 112350 2226 112378
rect 285166 112350 285194 112378
rect 98966 110110 98994 110138
rect 286006 109270 286034 109298
rect 2366 104958 2394 104986
rect 281750 104958 281778 104986
rect 281582 104902 281610 104930
rect 98910 103054 98938 103082
rect 3766 96110 3794 96138
rect 282646 96054 282674 96082
rect 292726 89558 292754 89586
rect 99022 88942 99050 88970
rect 98630 81886 98658 81914
rect 281918 76230 281946 76258
rect 2254 74942 2282 74970
rect 289366 69622 289394 69650
rect 99078 67774 99106 67802
rect 281974 63014 282002 63042
rect 98686 60718 98714 60746
rect 282030 56406 282058 56434
rect 2086 53718 2114 53746
rect 282086 49798 282114 49826
rect 98742 46606 98770 46634
rect 282142 43190 282170 43218
rect 98854 39550 98882 39578
rect 281806 36582 281834 36610
rect 2142 32606 2170 32634
rect 287686 29974 287714 30002
rect 2310 25550 2338 25578
rect 281862 23366 281890 23394
rect 98798 18382 98826 18410
rect 282198 16814 282226 16842
rect 2198 11438 2226 11466
rect 285166 10150 285194 10178
rect 2366 4382 2394 4410
rect 281750 3542 281778 3570
<< metal4 >>
rect -958 299086 -648 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 -648 299086
rect -958 299024 -648 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 -648 299024
rect -958 298962 -648 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 -648 298962
rect -958 298900 -648 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 -648 298900
rect -958 293175 -648 298872
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 -648 293175
rect -958 293113 -648 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 -648 293113
rect -958 293051 -648 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 -648 293051
rect -958 292989 -648 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 -648 292989
rect -958 284175 -648 292961
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 -648 284175
rect -958 284113 -648 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 -648 284113
rect -958 284051 -648 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 -648 284051
rect -958 283989 -648 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 -648 283989
rect -958 275175 -648 283961
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 -648 275175
rect -958 275113 -648 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 -648 275113
rect -958 275051 -648 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 -648 275051
rect -958 274989 -648 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 -648 274989
rect -958 266175 -648 274961
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 -648 266175
rect -958 266113 -648 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 -648 266113
rect -958 266051 -648 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 -648 266051
rect -958 265989 -648 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 -648 265989
rect -958 257175 -648 265961
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 -648 257175
rect -958 257113 -648 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 -648 257113
rect -958 257051 -648 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 -648 257051
rect -958 256989 -648 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 -648 256989
rect -958 248175 -648 256961
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 -648 248175
rect -958 248113 -648 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 -648 248113
rect -958 248051 -648 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 -648 248051
rect -958 247989 -648 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 -648 247989
rect -958 239175 -648 247961
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 -648 239175
rect -958 239113 -648 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 -648 239113
rect -958 239051 -648 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 -648 239051
rect -958 238989 -648 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 -648 238989
rect -958 230175 -648 238961
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 -648 230175
rect -958 230113 -648 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 -648 230113
rect -958 230051 -648 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 -648 230051
rect -958 229989 -648 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 -648 229989
rect -958 221175 -648 229961
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 -648 221175
rect -958 221113 -648 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 -648 221113
rect -958 221051 -648 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 -648 221051
rect -958 220989 -648 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 -648 220989
rect -958 212175 -648 220961
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 -648 212175
rect -958 212113 -648 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 -648 212113
rect -958 212051 -648 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 -648 212051
rect -958 211989 -648 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 -648 211989
rect -958 203175 -648 211961
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 -648 203175
rect -958 203113 -648 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 -648 203113
rect -958 203051 -648 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 -648 203051
rect -958 202989 -648 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 -648 202989
rect -958 194175 -648 202961
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 -648 194175
rect -958 194113 -648 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 -648 194113
rect -958 194051 -648 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 -648 194051
rect -958 193989 -648 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 -648 193989
rect -958 185175 -648 193961
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 -648 185175
rect -958 185113 -648 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 -648 185113
rect -958 185051 -648 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 -648 185051
rect -958 184989 -648 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 -648 184989
rect -958 176175 -648 184961
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 -648 176175
rect -958 176113 -648 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 -648 176113
rect -958 176051 -648 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 -648 176051
rect -958 175989 -648 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 -648 175989
rect -958 167175 -648 175961
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 -648 167175
rect -958 167113 -648 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 -648 167113
rect -958 167051 -648 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 -648 167051
rect -958 166989 -648 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 -648 166989
rect -958 158175 -648 166961
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 -648 158175
rect -958 158113 -648 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 -648 158113
rect -958 158051 -648 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 -648 158051
rect -958 157989 -648 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 -648 157989
rect -958 149175 -648 157961
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 -648 149175
rect -958 149113 -648 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 -648 149113
rect -958 149051 -648 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 -648 149051
rect -958 148989 -648 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 -648 148989
rect -958 140175 -648 148961
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 -648 140175
rect -958 140113 -648 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 -648 140113
rect -958 140051 -648 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 -648 140051
rect -958 139989 -648 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 -648 139989
rect -958 131175 -648 139961
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 -648 131175
rect -958 131113 -648 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 -648 131113
rect -958 131051 -648 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 -648 131051
rect -958 130989 -648 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 -648 130989
rect -958 122175 -648 130961
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 -648 122175
rect -958 122113 -648 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 -648 122113
rect -958 122051 -648 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 -648 122051
rect -958 121989 -648 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 -648 121989
rect -958 113175 -648 121961
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 -648 113175
rect -958 113113 -648 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 -648 113113
rect -958 113051 -648 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 -648 113051
rect -958 112989 -648 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 -648 112989
rect -958 104175 -648 112961
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 -648 104175
rect -958 104113 -648 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 -648 104113
rect -958 104051 -648 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 -648 104051
rect -958 103989 -648 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 -648 103989
rect -958 95175 -648 103961
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 -648 95175
rect -958 95113 -648 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 -648 95113
rect -958 95051 -648 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 -648 95051
rect -958 94989 -648 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 -648 94989
rect -958 86175 -648 94961
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 -648 86175
rect -958 86113 -648 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 -648 86113
rect -958 86051 -648 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 -648 86051
rect -958 85989 -648 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 -648 85989
rect -958 77175 -648 85961
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 -648 77175
rect -958 77113 -648 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 -648 77113
rect -958 77051 -648 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 -648 77051
rect -958 76989 -648 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 -648 76989
rect -958 68175 -648 76961
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 -648 68175
rect -958 68113 -648 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 -648 68113
rect -958 68051 -648 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 -648 68051
rect -958 67989 -648 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 -648 67989
rect -958 59175 -648 67961
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 -648 59175
rect -958 59113 -648 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 -648 59113
rect -958 59051 -648 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 -648 59051
rect -958 58989 -648 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 -648 58989
rect -958 50175 -648 58961
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 -648 50175
rect -958 50113 -648 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 -648 50113
rect -958 50051 -648 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 -648 50051
rect -958 49989 -648 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 -648 49989
rect -958 41175 -648 49961
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 -648 41175
rect -958 41113 -648 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 -648 41113
rect -958 41051 -648 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 -648 41051
rect -958 40989 -648 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 -648 40989
rect -958 32175 -648 40961
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 -648 32175
rect -958 32113 -648 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 -648 32113
rect -958 32051 -648 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 -648 32051
rect -958 31989 -648 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 -648 31989
rect -958 23175 -648 31961
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 -648 23175
rect -958 23113 -648 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 -648 23113
rect -958 23051 -648 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 -648 23051
rect -958 22989 -648 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 -648 22989
rect -958 14175 -648 22961
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 -648 14175
rect -958 14113 -648 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 -648 14113
rect -958 14051 -648 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 -648 14051
rect -958 13989 -648 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 -648 13989
rect -958 5175 -648 13961
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 -648 5175
rect -958 5113 -648 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 -648 5113
rect -958 5051 -648 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 -648 5051
rect -958 4989 -648 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 -648 4989
rect -958 -560 -648 4961
rect -478 298606 -168 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 -168 298606
rect -478 298544 -168 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 -168 298544
rect -478 298482 -168 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 -168 298482
rect -478 298420 -168 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 -168 298420
rect -478 290175 -168 298392
rect -478 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 -168 290175
rect -478 290113 -168 290147
rect -478 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 -168 290113
rect -478 290051 -168 290085
rect -478 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 -168 290051
rect -478 289989 -168 290023
rect -478 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 -168 289989
rect -478 281175 -168 289961
rect -478 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 -168 281175
rect -478 281113 -168 281147
rect -478 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 -168 281113
rect -478 281051 -168 281085
rect -478 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 -168 281051
rect -478 280989 -168 281023
rect -478 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 -168 280989
rect -478 272175 -168 280961
rect -478 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 -168 272175
rect -478 272113 -168 272147
rect -478 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 -168 272113
rect -478 272051 -168 272085
rect -478 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 -168 272051
rect -478 271989 -168 272023
rect -478 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 -168 271989
rect -478 263175 -168 271961
rect 2709 298606 3019 299134
rect 2709 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 3019 298606
rect 2709 298544 3019 298578
rect 2709 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 3019 298544
rect 2709 298482 3019 298516
rect 2709 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 3019 298482
rect 2709 298420 3019 298454
rect 2709 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 3019 298420
rect 2709 290175 3019 298392
rect 2709 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 3019 290175
rect 2709 290113 3019 290147
rect 2709 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 3019 290113
rect 2709 290051 3019 290085
rect 2709 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 3019 290051
rect 2709 289989 3019 290023
rect 2709 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 3019 289989
rect 2709 281175 3019 289961
rect 2709 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 3019 281175
rect 2709 281113 3019 281147
rect 2709 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 3019 281113
rect 2709 281051 3019 281085
rect 2709 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 3019 281051
rect 2709 280989 3019 281023
rect 2709 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 3019 280989
rect 2709 272175 3019 280961
rect 2709 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 3019 272175
rect 2709 272113 3019 272147
rect 2709 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 3019 272113
rect 2709 272051 3019 272085
rect 2709 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 3019 272051
rect 2709 271989 3019 272023
rect 2709 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 3019 271989
rect -478 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 -168 263175
rect -478 263113 -168 263147
rect -478 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 -168 263113
rect -478 263051 -168 263085
rect -478 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 -168 263051
rect -478 262989 -168 263023
rect -478 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 -168 262989
rect -478 254175 -168 262961
rect -478 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 -168 254175
rect -478 254113 -168 254147
rect -478 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 -168 254113
rect -478 254051 -168 254085
rect -478 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 -168 254051
rect -478 253989 -168 254023
rect -478 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 -168 253989
rect -478 245175 -168 253961
rect -478 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 -168 245175
rect -478 245113 -168 245147
rect -478 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 -168 245113
rect -478 245051 -168 245085
rect -478 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 -168 245051
rect -478 244989 -168 245023
rect -478 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 -168 244989
rect -478 236175 -168 244961
rect -478 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 -168 236175
rect -478 236113 -168 236147
rect -478 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 -168 236113
rect -478 236051 -168 236085
rect -478 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 -168 236051
rect -478 235989 -168 236023
rect -478 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 -168 235989
rect -478 227175 -168 235961
rect -478 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 -168 227175
rect -478 227113 -168 227147
rect -478 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 -168 227113
rect -478 227051 -168 227085
rect -478 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 -168 227051
rect -478 226989 -168 227023
rect -478 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 -168 226989
rect -478 218175 -168 226961
rect -478 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 -168 218175
rect -478 218113 -168 218147
rect -478 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 -168 218113
rect -478 218051 -168 218085
rect -478 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 -168 218051
rect -478 217989 -168 218023
rect -478 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 -168 217989
rect -478 209175 -168 217961
rect -478 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 -168 209175
rect -478 209113 -168 209147
rect -478 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 -168 209113
rect -478 209051 -168 209085
rect -478 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 -168 209051
rect -478 208989 -168 209023
rect -478 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 -168 208989
rect -478 200175 -168 208961
rect -478 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 -168 200175
rect -478 200113 -168 200147
rect -478 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 -168 200113
rect -478 200051 -168 200085
rect -478 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 -168 200051
rect -478 199989 -168 200023
rect -478 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 -168 199989
rect -478 191175 -168 199961
rect -478 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 -168 191175
rect -478 191113 -168 191147
rect -478 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 -168 191113
rect -478 191051 -168 191085
rect -478 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 -168 191051
rect -478 190989 -168 191023
rect -478 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 -168 190989
rect -478 182175 -168 190961
rect -478 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 -168 182175
rect -478 182113 -168 182147
rect -478 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 -168 182113
rect -478 182051 -168 182085
rect -478 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 -168 182051
rect -478 181989 -168 182023
rect -478 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 -168 181989
rect -478 173175 -168 181961
rect -478 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 -168 173175
rect -478 173113 -168 173147
rect -478 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 -168 173113
rect -478 173051 -168 173085
rect -478 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 -168 173051
rect -478 172989 -168 173023
rect -478 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 -168 172989
rect -478 164175 -168 172961
rect -478 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 -168 164175
rect -478 164113 -168 164147
rect -478 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 -168 164113
rect -478 164051 -168 164085
rect -478 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 -168 164051
rect -478 163989 -168 164023
rect -478 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 -168 163989
rect -478 155175 -168 163961
rect 2086 267610 2114 267615
rect 2086 159586 2114 267582
rect 2709 263175 3019 271961
rect 2709 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 3019 263175
rect 2709 263113 3019 263147
rect 2709 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 3019 263113
rect 2709 263051 3019 263085
rect 2709 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 3019 263051
rect 2709 262989 3019 263023
rect 2709 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 3019 262989
rect 2709 254175 3019 262961
rect 2709 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 3019 254175
rect 2709 254113 3019 254147
rect 2709 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 3019 254113
rect 2709 254051 3019 254085
rect 2709 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 3019 254051
rect 2709 253989 3019 254023
rect 2709 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 3019 253989
rect 2086 159553 2114 159558
rect 2142 245434 2170 245439
rect -478 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 -168 155175
rect -478 155113 -168 155147
rect -478 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 -168 155113
rect -478 155051 -168 155085
rect -478 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 -168 155051
rect -478 154989 -168 155023
rect -478 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 -168 154989
rect -478 146175 -168 154961
rect -478 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 -168 146175
rect -478 146113 -168 146147
rect -478 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 -168 146113
rect -478 146051 -168 146085
rect -478 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 -168 146051
rect -478 145989 -168 146023
rect -478 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 -168 145989
rect -478 137175 -168 145961
rect -478 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 -168 137175
rect -478 137113 -168 137147
rect -478 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 -168 137113
rect -478 137051 -168 137085
rect -478 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 -168 137051
rect -478 136989 -168 137023
rect -478 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 -168 136989
rect -478 128175 -168 136961
rect -478 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 -168 128175
rect -478 128113 -168 128147
rect -478 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 -168 128113
rect -478 128051 -168 128085
rect -478 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 -168 128051
rect -478 127989 -168 128023
rect -478 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 -168 127989
rect -478 119175 -168 127961
rect -478 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 -168 119175
rect -478 119113 -168 119147
rect -478 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 -168 119113
rect -478 119051 -168 119085
rect -478 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 -168 119051
rect -478 118989 -168 119023
rect -478 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 -168 118989
rect -478 110175 -168 118961
rect -478 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 -168 110175
rect -478 110113 -168 110147
rect -478 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 -168 110113
rect -478 110051 -168 110085
rect -478 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 -168 110051
rect -478 109989 -168 110023
rect -478 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 -168 109989
rect -478 101175 -168 109961
rect -478 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 -168 101175
rect -478 101113 -168 101147
rect -478 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 -168 101113
rect -478 101051 -168 101085
rect -478 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 -168 101051
rect -478 100989 -168 101023
rect -478 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 -168 100989
rect -478 92175 -168 100961
rect -478 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 -168 92175
rect -478 92113 -168 92147
rect -478 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 -168 92113
rect -478 92051 -168 92085
rect -478 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 -168 92051
rect -478 91989 -168 92023
rect -478 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 -168 91989
rect -478 83175 -168 91961
rect -478 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 -168 83175
rect -478 83113 -168 83147
rect -478 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 -168 83113
rect -478 83051 -168 83085
rect -478 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 -168 83051
rect -478 82989 -168 83023
rect -478 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 -168 82989
rect -478 74175 -168 82961
rect -478 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 -168 74175
rect -478 74113 -168 74147
rect -478 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 -168 74113
rect -478 74051 -168 74085
rect -478 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 -168 74051
rect -478 73989 -168 74023
rect -478 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 -168 73989
rect -478 65175 -168 73961
rect -478 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 -168 65175
rect -478 65113 -168 65147
rect -478 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 -168 65113
rect -478 65051 -168 65085
rect -478 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 -168 65051
rect -478 64989 -168 65023
rect -478 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 -168 64989
rect -478 56175 -168 64961
rect -478 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 -168 56175
rect -478 56113 -168 56147
rect -478 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 -168 56113
rect -478 56051 -168 56085
rect -478 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 -168 56051
rect -478 55989 -168 56023
rect -478 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 -168 55989
rect -478 47175 -168 55961
rect 2086 156730 2114 156735
rect 2086 53746 2114 156702
rect 2142 138474 2170 245406
rect 2709 245175 3019 253961
rect 2709 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 3019 245175
rect 2709 245113 3019 245147
rect 2709 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 3019 245113
rect 2709 245051 3019 245085
rect 2709 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 3019 245051
rect 2709 244989 3019 245023
rect 2709 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 3019 244989
rect 2709 236175 3019 244961
rect 2709 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 3019 236175
rect 2709 236113 3019 236147
rect 2709 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 3019 236113
rect 2709 236051 3019 236085
rect 2709 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 3019 236051
rect 2709 235989 3019 236023
rect 2709 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 3019 235989
rect 2709 227175 3019 235961
rect 2709 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 3019 227175
rect 2709 227113 3019 227147
rect 2709 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 3019 227113
rect 2709 227051 3019 227085
rect 2709 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 3019 227051
rect 2709 226989 3019 227023
rect 2709 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 3019 226989
rect 2142 138441 2170 138446
rect 2198 223258 2226 223263
rect 2086 53713 2114 53718
rect 2142 134554 2170 134559
rect -478 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 -168 47175
rect -478 47113 -168 47147
rect -478 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 -168 47113
rect -478 47051 -168 47085
rect -478 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 -168 47051
rect -478 46989 -168 47023
rect -478 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 -168 46989
rect -478 38175 -168 46961
rect -478 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 -168 38175
rect -478 38113 -168 38147
rect -478 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 -168 38113
rect -478 38051 -168 38085
rect -478 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 -168 38051
rect -478 37989 -168 38023
rect -478 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 -168 37989
rect -478 29175 -168 37961
rect 2142 32634 2170 134526
rect 2198 117306 2226 223230
rect 2709 218175 3019 226961
rect 2709 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 3019 218175
rect 2709 218113 3019 218147
rect 2709 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 3019 218113
rect 2709 218051 3019 218085
rect 2709 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 3019 218051
rect 2709 217989 3019 218023
rect 2709 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 3019 217989
rect 2709 209175 3019 217961
rect 2709 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 3019 209175
rect 2709 209113 3019 209147
rect 2709 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 3019 209113
rect 2709 209051 3019 209085
rect 2709 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 3019 209051
rect 2709 208989 3019 209023
rect 2709 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 3019 208989
rect 2709 200175 3019 208961
rect 4569 299086 4879 299134
rect 4569 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 4879 299086
rect 4569 299024 4879 299058
rect 4569 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 4879 299024
rect 4569 298962 4879 298996
rect 4569 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 4879 298962
rect 4569 298900 4879 298934
rect 4569 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 4879 298900
rect 4569 293175 4879 298872
rect 4569 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 4879 293175
rect 4569 293113 4879 293147
rect 4569 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 4879 293113
rect 4569 293051 4879 293085
rect 4569 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 4879 293051
rect 4569 292989 4879 293023
rect 4569 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 4879 292989
rect 4569 284175 4879 292961
rect 4569 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 4879 284175
rect 4569 284113 4879 284147
rect 4569 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 4879 284113
rect 4569 284051 4879 284085
rect 4569 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 4879 284051
rect 4569 283989 4879 284023
rect 4569 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 4879 283989
rect 4569 275175 4879 283961
rect 4569 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 4879 275175
rect 4569 275113 4879 275147
rect 4569 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 4879 275113
rect 4569 275051 4879 275085
rect 4569 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 4879 275051
rect 4569 274989 4879 275023
rect 4569 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 4879 274989
rect 4569 266175 4879 274961
rect 4569 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 4879 266175
rect 4569 266113 4879 266147
rect 4569 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 4879 266113
rect 4569 266051 4879 266085
rect 4569 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 4879 266051
rect 4569 265989 4879 266023
rect 4569 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 4879 265989
rect 4569 257175 4879 265961
rect 4569 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 4879 257175
rect 4569 257113 4879 257147
rect 4569 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 4879 257113
rect 4569 257051 4879 257085
rect 4569 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 4879 257051
rect 4569 256989 4879 257023
rect 4569 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 4879 256989
rect 4569 248175 4879 256961
rect 4569 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 4879 248175
rect 4569 248113 4879 248147
rect 4569 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 4879 248113
rect 4569 248051 4879 248085
rect 4569 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 4879 248051
rect 4569 247989 4879 248023
rect 4569 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 4879 247989
rect 4569 239175 4879 247961
rect 4569 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 4879 239175
rect 4569 239113 4879 239147
rect 4569 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 4879 239113
rect 4569 239051 4879 239085
rect 4569 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 4879 239051
rect 4569 238989 4879 239023
rect 4569 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 4879 238989
rect 4569 230175 4879 238961
rect 4569 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 4879 230175
rect 4569 230113 4879 230147
rect 4569 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 4879 230113
rect 4569 230051 4879 230085
rect 4569 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 4879 230051
rect 4569 229989 4879 230023
rect 4569 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 4879 229989
rect 4569 221175 4879 229961
rect 4569 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 4879 221175
rect 4569 221113 4879 221147
rect 4569 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 4879 221113
rect 4569 221051 4879 221085
rect 4569 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 4879 221051
rect 4569 220989 4879 221023
rect 4569 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 4879 220989
rect 4569 212175 4879 220961
rect 4569 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 4879 212175
rect 4569 212113 4879 212147
rect 4569 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 4879 212113
rect 4569 212051 4879 212085
rect 4569 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 4879 212051
rect 4569 211989 4879 212023
rect 4569 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 4879 211989
rect 4569 203175 4879 211961
rect 4569 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 4879 203175
rect 4569 203113 4879 203147
rect 4569 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 4879 203113
rect 4569 203051 4879 203085
rect 4569 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 4879 203051
rect 4569 202989 4879 203023
rect 4569 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 4879 202989
rect 2709 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 3019 200175
rect 2709 200113 3019 200147
rect 2709 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 3019 200113
rect 2709 200051 3019 200085
rect 2709 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 3019 200051
rect 2709 199989 3019 200023
rect 2709 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 3019 199989
rect 2709 191175 3019 199961
rect 2709 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 3019 191175
rect 2709 191113 3019 191147
rect 2709 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 3019 191113
rect 2709 191051 3019 191085
rect 2709 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 3019 191051
rect 2709 190989 3019 191023
rect 2709 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 3019 190989
rect 2709 182175 3019 190961
rect 2709 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 3019 182175
rect 2709 182113 3019 182147
rect 2709 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 3019 182113
rect 2709 182051 3019 182085
rect 2709 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 3019 182051
rect 2709 181989 3019 182023
rect 2709 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 3019 181989
rect 2198 117273 2226 117278
rect 2254 178906 2282 178911
rect 2142 32601 2170 32606
rect 2198 112378 2226 112383
rect -478 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 -168 29175
rect -478 29113 -168 29147
rect -478 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 -168 29113
rect -478 29051 -168 29085
rect -478 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 -168 29051
rect -478 28989 -168 29023
rect -478 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 -168 28989
rect -478 20175 -168 28961
rect -478 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 -168 20175
rect -478 20113 -168 20147
rect -478 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 -168 20113
rect -478 20051 -168 20085
rect -478 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 -168 20051
rect -478 19989 -168 20023
rect -478 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 -168 19989
rect -478 11175 -168 19961
rect 2198 11466 2226 112350
rect 2254 74970 2282 178878
rect 2709 173175 3019 181961
rect 2709 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 3019 173175
rect 2709 173113 3019 173147
rect 2709 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 3019 173113
rect 2709 173051 3019 173085
rect 2709 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 3019 173051
rect 2709 172989 3019 173023
rect 2709 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 3019 172989
rect 2709 164175 3019 172961
rect 2709 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 3019 164175
rect 2709 164113 3019 164147
rect 2709 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 3019 164113
rect 2709 164051 3019 164085
rect 2709 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 3019 164051
rect 2709 163989 3019 164023
rect 2709 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 3019 163989
rect 2709 155175 3019 163961
rect 2709 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 3019 155175
rect 2709 155113 3019 155147
rect 2709 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 3019 155113
rect 2709 155051 3019 155085
rect 2709 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 3019 155051
rect 2709 154989 3019 155023
rect 2709 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 3019 154989
rect 2709 146175 3019 154961
rect 2709 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 3019 146175
rect 2709 146113 3019 146147
rect 2709 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 3019 146113
rect 2709 146051 3019 146085
rect 2709 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 3019 146051
rect 2709 145989 3019 146023
rect 2709 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 3019 145989
rect 2709 137175 3019 145961
rect 2709 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 3019 137175
rect 2709 137113 3019 137147
rect 2709 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 3019 137113
rect 2709 137051 3019 137085
rect 2709 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 3019 137051
rect 2709 136989 3019 137023
rect 2709 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 3019 136989
rect 2709 128175 3019 136961
rect 2709 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 3019 128175
rect 2709 128113 3019 128147
rect 2709 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 3019 128113
rect 2709 128051 3019 128085
rect 2709 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 3019 128051
rect 2709 127989 3019 128023
rect 2709 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 3019 127989
rect 2254 74937 2282 74942
rect 2310 127162 2338 127167
rect 2310 25578 2338 127134
rect 2709 119175 3019 127961
rect 2709 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 3019 119175
rect 2709 119113 3019 119147
rect 2709 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 3019 119113
rect 2709 119051 3019 119085
rect 2709 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 3019 119051
rect 2709 118989 3019 119023
rect 2709 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 3019 118989
rect 2709 110175 3019 118961
rect 2709 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 3019 110175
rect 2709 110113 3019 110147
rect 2709 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 3019 110113
rect 2709 110051 3019 110085
rect 2709 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 3019 110051
rect 2709 109989 3019 110023
rect 2709 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 3019 109989
rect 2310 25545 2338 25550
rect 2366 104986 2394 104991
rect 2198 11433 2226 11438
rect -478 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 -168 11175
rect -478 11113 -168 11147
rect -478 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 -168 11113
rect -478 11051 -168 11085
rect -478 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 -168 11051
rect -478 10989 -168 11023
rect -478 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 -168 10989
rect -478 2175 -168 10961
rect 2366 4410 2394 104958
rect 2366 4377 2394 4382
rect 2709 101175 3019 109961
rect 2709 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 3019 101175
rect 2709 101113 3019 101147
rect 2709 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 3019 101113
rect 2709 101051 3019 101085
rect 2709 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 3019 101051
rect 2709 100989 3019 101023
rect 2709 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 3019 100989
rect 2709 92175 3019 100961
rect 3766 201082 3794 201087
rect 3766 96138 3794 201054
rect 3766 96105 3794 96110
rect 4569 194175 4879 202961
rect 4569 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 4879 194175
rect 4569 194113 4879 194147
rect 4569 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 4879 194113
rect 4569 194051 4879 194085
rect 4569 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 4879 194051
rect 4569 193989 4879 194023
rect 4569 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 4879 193989
rect 4569 185175 4879 193961
rect 4569 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 4879 185175
rect 4569 185113 4879 185147
rect 4569 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 4879 185113
rect 4569 185051 4879 185085
rect 4569 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 4879 185051
rect 4569 184989 4879 185023
rect 4569 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 4879 184989
rect 4569 176175 4879 184961
rect 4569 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 4879 176175
rect 4569 176113 4879 176147
rect 4569 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 4879 176113
rect 4569 176051 4879 176085
rect 4569 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 4879 176051
rect 4569 175989 4879 176023
rect 4569 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 4879 175989
rect 4569 167175 4879 175961
rect 4569 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 4879 167175
rect 4569 167113 4879 167147
rect 4569 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 4879 167113
rect 4569 167051 4879 167085
rect 4569 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 4879 167051
rect 4569 166989 4879 167023
rect 4569 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 4879 166989
rect 4569 158175 4879 166961
rect 4569 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 4879 158175
rect 4569 158113 4879 158147
rect 4569 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 4879 158113
rect 4569 158051 4879 158085
rect 4569 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 4879 158051
rect 4569 157989 4879 158023
rect 4569 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 4879 157989
rect 4569 149175 4879 157961
rect 4569 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 4879 149175
rect 4569 149113 4879 149147
rect 4569 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 4879 149113
rect 4569 149051 4879 149085
rect 4569 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 4879 149051
rect 4569 148989 4879 149023
rect 4569 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 4879 148989
rect 4569 140175 4879 148961
rect 4569 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 4879 140175
rect 4569 140113 4879 140147
rect 4569 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 4879 140113
rect 4569 140051 4879 140085
rect 4569 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 4879 140051
rect 4569 139989 4879 140023
rect 4569 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 4879 139989
rect 4569 131175 4879 139961
rect 4569 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 4879 131175
rect 4569 131113 4879 131147
rect 4569 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 4879 131113
rect 4569 131051 4879 131085
rect 4569 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 4879 131051
rect 4569 130989 4879 131023
rect 4569 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 4879 130989
rect 4569 122175 4879 130961
rect 4569 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 4879 122175
rect 4569 122113 4879 122147
rect 4569 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 4879 122113
rect 4569 122051 4879 122085
rect 4569 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 4879 122051
rect 4569 121989 4879 122023
rect 4569 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 4879 121989
rect 4569 113175 4879 121961
rect 4569 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 4879 113175
rect 4569 113113 4879 113147
rect 4569 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 4879 113113
rect 4569 113051 4879 113085
rect 4569 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 4879 113051
rect 4569 112989 4879 113023
rect 4569 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 4879 112989
rect 4569 104175 4879 112961
rect 4569 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 4879 104175
rect 4569 104113 4879 104147
rect 4569 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 4879 104113
rect 4569 104051 4879 104085
rect 4569 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 4879 104051
rect 4569 103989 4879 104023
rect 4569 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 4879 103989
rect 2709 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 3019 92175
rect 2709 92113 3019 92147
rect 2709 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 3019 92113
rect 2709 92051 3019 92085
rect 2709 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 3019 92051
rect 2709 91989 3019 92023
rect 2709 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 3019 91989
rect 2709 83175 3019 91961
rect 2709 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 3019 83175
rect 2709 83113 3019 83147
rect 2709 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 3019 83113
rect 2709 83051 3019 83085
rect 2709 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 3019 83051
rect 2709 82989 3019 83023
rect 2709 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 3019 82989
rect 2709 74175 3019 82961
rect 2709 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 3019 74175
rect 2709 74113 3019 74147
rect 2709 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 3019 74113
rect 2709 74051 3019 74085
rect 2709 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 3019 74051
rect 2709 73989 3019 74023
rect 2709 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 3019 73989
rect 2709 65175 3019 73961
rect 2709 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 3019 65175
rect 2709 65113 3019 65147
rect 2709 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 3019 65113
rect 2709 65051 3019 65085
rect 2709 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 3019 65051
rect 2709 64989 3019 65023
rect 2709 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 3019 64989
rect 2709 56175 3019 64961
rect 2709 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 3019 56175
rect 2709 56113 3019 56147
rect 2709 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 3019 56113
rect 2709 56051 3019 56085
rect 2709 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 3019 56051
rect 2709 55989 3019 56023
rect 2709 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 3019 55989
rect 2709 47175 3019 55961
rect 2709 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 3019 47175
rect 2709 47113 3019 47147
rect 2709 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 3019 47113
rect 2709 47051 3019 47085
rect 2709 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 3019 47051
rect 2709 46989 3019 47023
rect 2709 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 3019 46989
rect 2709 38175 3019 46961
rect 2709 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 3019 38175
rect 2709 38113 3019 38147
rect 2709 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 3019 38113
rect 2709 38051 3019 38085
rect 2709 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 3019 38051
rect 2709 37989 3019 38023
rect 2709 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 3019 37989
rect 2709 29175 3019 37961
rect 2709 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 3019 29175
rect 2709 29113 3019 29147
rect 2709 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 3019 29113
rect 2709 29051 3019 29085
rect 2709 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 3019 29051
rect 2709 28989 3019 29023
rect 2709 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 3019 28989
rect 2709 20175 3019 28961
rect 2709 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 3019 20175
rect 2709 20113 3019 20147
rect 2709 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 3019 20113
rect 2709 20051 3019 20085
rect 2709 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 3019 20051
rect 2709 19989 3019 20023
rect 2709 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 3019 19989
rect 2709 11175 3019 19961
rect 2709 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 3019 11175
rect 2709 11113 3019 11147
rect 2709 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 3019 11113
rect 2709 11051 3019 11085
rect 2709 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 3019 11051
rect 2709 10989 3019 11023
rect 2709 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 3019 10989
rect -478 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 -168 2175
rect -478 2113 -168 2147
rect -478 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 -168 2113
rect -478 2051 -168 2085
rect -478 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 -168 2051
rect -478 1989 -168 2023
rect -478 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 -168 1989
rect -478 -80 -168 1961
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 -168 -80
rect -478 -142 -168 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 -168 -142
rect -478 -204 -168 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 -168 -204
rect -478 -266 -168 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 -168 -266
rect -478 -342 -168 -294
rect 2709 2175 3019 10961
rect 2709 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 3019 2175
rect 2709 2113 3019 2147
rect 2709 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 3019 2113
rect 2709 2051 3019 2085
rect 2709 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 3019 2051
rect 2709 1989 3019 2023
rect 2709 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 3019 1989
rect 2709 -80 3019 1961
rect 2709 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 3019 -80
rect 2709 -142 3019 -108
rect 2709 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 3019 -142
rect 2709 -204 3019 -170
rect 2709 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 3019 -204
rect 2709 -266 3019 -232
rect 2709 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 3019 -266
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 -648 -560
rect -958 -622 -648 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 -648 -622
rect -958 -684 -648 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 -648 -684
rect -958 -746 -648 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 -648 -746
rect -958 -822 -648 -774
rect 2709 -822 3019 -294
rect 4569 95175 4879 103961
rect 4569 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 4879 95175
rect 4569 95113 4879 95147
rect 4569 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 4879 95113
rect 4569 95051 4879 95085
rect 4569 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 4879 95051
rect 4569 94989 4879 95023
rect 4569 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 4879 94989
rect 4569 86175 4879 94961
rect 4569 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 4879 86175
rect 4569 86113 4879 86147
rect 4569 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 4879 86113
rect 4569 86051 4879 86085
rect 4569 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 4879 86051
rect 4569 85989 4879 86023
rect 4569 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 4879 85989
rect 4569 77175 4879 85961
rect 4569 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 4879 77175
rect 4569 77113 4879 77147
rect 4569 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 4879 77113
rect 4569 77051 4879 77085
rect 4569 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 4879 77051
rect 4569 76989 4879 77023
rect 4569 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 4879 76989
rect 4569 68175 4879 76961
rect 4569 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 4879 68175
rect 4569 68113 4879 68147
rect 4569 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 4879 68113
rect 4569 68051 4879 68085
rect 4569 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 4879 68051
rect 4569 67989 4879 68023
rect 4569 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 4879 67989
rect 4569 59175 4879 67961
rect 4569 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 4879 59175
rect 4569 59113 4879 59147
rect 4569 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 4879 59113
rect 4569 59051 4879 59085
rect 4569 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 4879 59051
rect 4569 58989 4879 59023
rect 4569 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 4879 58989
rect 4569 50175 4879 58961
rect 4569 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 4879 50175
rect 4569 50113 4879 50147
rect 4569 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 4879 50113
rect 4569 50051 4879 50085
rect 4569 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 4879 50051
rect 4569 49989 4879 50023
rect 4569 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 4879 49989
rect 4569 41175 4879 49961
rect 4569 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 4879 41175
rect 4569 41113 4879 41147
rect 4569 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 4879 41113
rect 4569 41051 4879 41085
rect 4569 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 4879 41051
rect 4569 40989 4879 41023
rect 4569 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 4879 40989
rect 4569 32175 4879 40961
rect 4569 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 4879 32175
rect 4569 32113 4879 32147
rect 4569 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 4879 32113
rect 4569 32051 4879 32085
rect 4569 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 4879 32051
rect 4569 31989 4879 32023
rect 4569 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 4879 31989
rect 4569 23175 4879 31961
rect 4569 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 4879 23175
rect 4569 23113 4879 23147
rect 4569 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 4879 23113
rect 4569 23051 4879 23085
rect 4569 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 4879 23051
rect 4569 22989 4879 23023
rect 4569 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 4879 22989
rect 4569 14175 4879 22961
rect 4569 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 4879 14175
rect 4569 14113 4879 14147
rect 4569 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 4879 14113
rect 4569 14051 4879 14085
rect 4569 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 4879 14051
rect 4569 13989 4879 14023
rect 4569 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 4879 13989
rect 4569 5175 4879 13961
rect 4569 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 4879 5175
rect 4569 5113 4879 5147
rect 4569 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 4879 5113
rect 4569 5051 4879 5085
rect 4569 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 4879 5051
rect 4569 4989 4879 5023
rect 4569 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 4879 4989
rect 4569 -560 4879 4961
rect 4569 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 4879 -560
rect 4569 -622 4879 -588
rect 4569 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 4879 -622
rect 4569 -684 4879 -650
rect 4569 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 4879 -684
rect 4569 -746 4879 -712
rect 4569 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 4879 -746
rect 4569 -822 4879 -774
rect 18069 298606 18379 299134
rect 18069 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 18379 298606
rect 18069 298544 18379 298578
rect 18069 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 18379 298544
rect 18069 298482 18379 298516
rect 18069 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 18379 298482
rect 18069 298420 18379 298454
rect 18069 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 18379 298420
rect 18069 290175 18379 298392
rect 18069 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 18379 290175
rect 18069 290113 18379 290147
rect 18069 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 18379 290113
rect 18069 290051 18379 290085
rect 18069 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 18379 290051
rect 18069 289989 18379 290023
rect 18069 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 18379 289989
rect 18069 281175 18379 289961
rect 18069 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 18379 281175
rect 18069 281113 18379 281147
rect 18069 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 18379 281113
rect 18069 281051 18379 281085
rect 18069 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 18379 281051
rect 18069 280989 18379 281023
rect 18069 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 18379 280989
rect 18069 272175 18379 280961
rect 18069 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 18379 272175
rect 18069 272113 18379 272147
rect 18069 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 18379 272113
rect 18069 272051 18379 272085
rect 18069 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 18379 272051
rect 18069 271989 18379 272023
rect 18069 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 18379 271989
rect 18069 263175 18379 271961
rect 18069 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 18379 263175
rect 18069 263113 18379 263147
rect 18069 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 18379 263113
rect 18069 263051 18379 263085
rect 18069 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 18379 263051
rect 18069 262989 18379 263023
rect 18069 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 18379 262989
rect 18069 254175 18379 262961
rect 18069 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 18379 254175
rect 18069 254113 18379 254147
rect 18069 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 18379 254113
rect 18069 254051 18379 254085
rect 18069 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 18379 254051
rect 18069 253989 18379 254023
rect 18069 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 18379 253989
rect 18069 245175 18379 253961
rect 18069 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 18379 245175
rect 18069 245113 18379 245147
rect 18069 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 18379 245113
rect 18069 245051 18379 245085
rect 18069 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 18379 245051
rect 18069 244989 18379 245023
rect 18069 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 18379 244989
rect 18069 236175 18379 244961
rect 18069 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 18379 236175
rect 18069 236113 18379 236147
rect 18069 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 18379 236113
rect 18069 236051 18379 236085
rect 18069 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 18379 236051
rect 18069 235989 18379 236023
rect 18069 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 18379 235989
rect 18069 227175 18379 235961
rect 18069 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 18379 227175
rect 18069 227113 18379 227147
rect 18069 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 18379 227113
rect 18069 227051 18379 227085
rect 18069 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 18379 227051
rect 18069 226989 18379 227023
rect 18069 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 18379 226989
rect 18069 218175 18379 226961
rect 18069 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 18379 218175
rect 18069 218113 18379 218147
rect 18069 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 18379 218113
rect 18069 218051 18379 218085
rect 18069 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 18379 218051
rect 18069 217989 18379 218023
rect 18069 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 18379 217989
rect 18069 209175 18379 217961
rect 18069 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 18379 209175
rect 18069 209113 18379 209147
rect 18069 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 18379 209113
rect 18069 209051 18379 209085
rect 18069 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 18379 209051
rect 18069 208989 18379 209023
rect 18069 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 18379 208989
rect 18069 200175 18379 208961
rect 18069 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 18379 200175
rect 18069 200113 18379 200147
rect 18069 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 18379 200113
rect 18069 200051 18379 200085
rect 18069 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 18379 200051
rect 18069 199989 18379 200023
rect 18069 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 18379 199989
rect 18069 191175 18379 199961
rect 18069 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 18379 191175
rect 18069 191113 18379 191147
rect 18069 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 18379 191113
rect 18069 191051 18379 191085
rect 18069 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 18379 191051
rect 18069 190989 18379 191023
rect 18069 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 18379 190989
rect 18069 182175 18379 190961
rect 18069 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 18379 182175
rect 18069 182113 18379 182147
rect 18069 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 18379 182113
rect 18069 182051 18379 182085
rect 18069 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 18379 182051
rect 18069 181989 18379 182023
rect 18069 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 18379 181989
rect 18069 173175 18379 181961
rect 18069 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 18379 173175
rect 18069 173113 18379 173147
rect 18069 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 18379 173113
rect 18069 173051 18379 173085
rect 18069 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 18379 173051
rect 18069 172989 18379 173023
rect 18069 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 18379 172989
rect 18069 164175 18379 172961
rect 18069 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 18379 164175
rect 18069 164113 18379 164147
rect 18069 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 18379 164113
rect 18069 164051 18379 164085
rect 18069 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 18379 164051
rect 18069 163989 18379 164023
rect 18069 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 18379 163989
rect 18069 155175 18379 163961
rect 18069 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 18379 155175
rect 18069 155113 18379 155147
rect 18069 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 18379 155113
rect 18069 155051 18379 155085
rect 18069 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 18379 155051
rect 18069 154989 18379 155023
rect 18069 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 18379 154989
rect 18069 146175 18379 154961
rect 18069 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 18379 146175
rect 18069 146113 18379 146147
rect 18069 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 18379 146113
rect 18069 146051 18379 146085
rect 18069 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 18379 146051
rect 18069 145989 18379 146023
rect 18069 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 18379 145989
rect 18069 137175 18379 145961
rect 18069 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 18379 137175
rect 18069 137113 18379 137147
rect 18069 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 18379 137113
rect 18069 137051 18379 137085
rect 18069 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 18379 137051
rect 18069 136989 18379 137023
rect 18069 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 18379 136989
rect 18069 128175 18379 136961
rect 18069 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 18379 128175
rect 18069 128113 18379 128147
rect 18069 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 18379 128113
rect 18069 128051 18379 128085
rect 18069 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 18379 128051
rect 18069 127989 18379 128023
rect 18069 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 18379 127989
rect 18069 119175 18379 127961
rect 18069 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 18379 119175
rect 18069 119113 18379 119147
rect 18069 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 18379 119113
rect 18069 119051 18379 119085
rect 18069 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 18379 119051
rect 18069 118989 18379 119023
rect 18069 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 18379 118989
rect 18069 110175 18379 118961
rect 18069 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 18379 110175
rect 18069 110113 18379 110147
rect 18069 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 18379 110113
rect 18069 110051 18379 110085
rect 18069 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 18379 110051
rect 18069 109989 18379 110023
rect 18069 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 18379 109989
rect 18069 101175 18379 109961
rect 18069 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 18379 101175
rect 18069 101113 18379 101147
rect 18069 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 18379 101113
rect 18069 101051 18379 101085
rect 18069 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 18379 101051
rect 18069 100989 18379 101023
rect 18069 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 18379 100989
rect 18069 92175 18379 100961
rect 18069 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 18379 92175
rect 18069 92113 18379 92147
rect 18069 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 18379 92113
rect 18069 92051 18379 92085
rect 18069 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 18379 92051
rect 18069 91989 18379 92023
rect 18069 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 18379 91989
rect 18069 83175 18379 91961
rect 18069 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 18379 83175
rect 18069 83113 18379 83147
rect 18069 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 18379 83113
rect 18069 83051 18379 83085
rect 18069 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 18379 83051
rect 18069 82989 18379 83023
rect 18069 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 18379 82989
rect 18069 74175 18379 82961
rect 18069 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 18379 74175
rect 18069 74113 18379 74147
rect 18069 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 18379 74113
rect 18069 74051 18379 74085
rect 18069 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 18379 74051
rect 18069 73989 18379 74023
rect 18069 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 18379 73989
rect 18069 65175 18379 73961
rect 18069 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 18379 65175
rect 18069 65113 18379 65147
rect 18069 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 18379 65113
rect 18069 65051 18379 65085
rect 18069 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 18379 65051
rect 18069 64989 18379 65023
rect 18069 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 18379 64989
rect 18069 56175 18379 64961
rect 18069 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 18379 56175
rect 18069 56113 18379 56147
rect 18069 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 18379 56113
rect 18069 56051 18379 56085
rect 18069 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 18379 56051
rect 18069 55989 18379 56023
rect 18069 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 18379 55989
rect 18069 47175 18379 55961
rect 18069 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 18379 47175
rect 18069 47113 18379 47147
rect 18069 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 18379 47113
rect 18069 47051 18379 47085
rect 18069 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 18379 47051
rect 18069 46989 18379 47023
rect 18069 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 18379 46989
rect 18069 38175 18379 46961
rect 18069 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 18379 38175
rect 18069 38113 18379 38147
rect 18069 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 18379 38113
rect 18069 38051 18379 38085
rect 18069 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 18379 38051
rect 18069 37989 18379 38023
rect 18069 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 18379 37989
rect 18069 29175 18379 37961
rect 18069 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 18379 29175
rect 18069 29113 18379 29147
rect 18069 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 18379 29113
rect 18069 29051 18379 29085
rect 18069 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 18379 29051
rect 18069 28989 18379 29023
rect 18069 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 18379 28989
rect 18069 20175 18379 28961
rect 18069 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 18379 20175
rect 18069 20113 18379 20147
rect 18069 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 18379 20113
rect 18069 20051 18379 20085
rect 18069 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 18379 20051
rect 18069 19989 18379 20023
rect 18069 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 18379 19989
rect 18069 11175 18379 19961
rect 18069 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 18379 11175
rect 18069 11113 18379 11147
rect 18069 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 18379 11113
rect 18069 11051 18379 11085
rect 18069 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 18379 11051
rect 18069 10989 18379 11023
rect 18069 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 18379 10989
rect 18069 2175 18379 10961
rect 18069 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 18379 2175
rect 18069 2113 18379 2147
rect 18069 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 18379 2113
rect 18069 2051 18379 2085
rect 18069 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 18379 2051
rect 18069 1989 18379 2023
rect 18069 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 18379 1989
rect 18069 -80 18379 1961
rect 18069 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 18379 -80
rect 18069 -142 18379 -108
rect 18069 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 18379 -142
rect 18069 -204 18379 -170
rect 18069 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 18379 -204
rect 18069 -266 18379 -232
rect 18069 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 18379 -266
rect 18069 -822 18379 -294
rect 19929 299086 20239 299134
rect 19929 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 20239 299086
rect 19929 299024 20239 299058
rect 19929 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 20239 299024
rect 19929 298962 20239 298996
rect 19929 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 20239 298962
rect 19929 298900 20239 298934
rect 19929 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 20239 298900
rect 19929 293175 20239 298872
rect 19929 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 20239 293175
rect 19929 293113 20239 293147
rect 19929 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 20239 293113
rect 19929 293051 20239 293085
rect 19929 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 20239 293051
rect 19929 292989 20239 293023
rect 19929 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 20239 292989
rect 19929 284175 20239 292961
rect 19929 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 20239 284175
rect 19929 284113 20239 284147
rect 19929 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 20239 284113
rect 19929 284051 20239 284085
rect 19929 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 20239 284051
rect 19929 283989 20239 284023
rect 19929 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 20239 283989
rect 19929 275175 20239 283961
rect 19929 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 20239 275175
rect 19929 275113 20239 275147
rect 19929 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 20239 275113
rect 19929 275051 20239 275085
rect 19929 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 20239 275051
rect 19929 274989 20239 275023
rect 19929 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 20239 274989
rect 19929 266175 20239 274961
rect 19929 266147 19977 266175
rect 20005 266147 20039 266175
rect 20067 266147 20101 266175
rect 20129 266147 20163 266175
rect 20191 266147 20239 266175
rect 19929 266113 20239 266147
rect 19929 266085 19977 266113
rect 20005 266085 20039 266113
rect 20067 266085 20101 266113
rect 20129 266085 20163 266113
rect 20191 266085 20239 266113
rect 19929 266051 20239 266085
rect 19929 266023 19977 266051
rect 20005 266023 20039 266051
rect 20067 266023 20101 266051
rect 20129 266023 20163 266051
rect 20191 266023 20239 266051
rect 19929 265989 20239 266023
rect 19929 265961 19977 265989
rect 20005 265961 20039 265989
rect 20067 265961 20101 265989
rect 20129 265961 20163 265989
rect 20191 265961 20239 265989
rect 19929 257175 20239 265961
rect 19929 257147 19977 257175
rect 20005 257147 20039 257175
rect 20067 257147 20101 257175
rect 20129 257147 20163 257175
rect 20191 257147 20239 257175
rect 19929 257113 20239 257147
rect 19929 257085 19977 257113
rect 20005 257085 20039 257113
rect 20067 257085 20101 257113
rect 20129 257085 20163 257113
rect 20191 257085 20239 257113
rect 19929 257051 20239 257085
rect 19929 257023 19977 257051
rect 20005 257023 20039 257051
rect 20067 257023 20101 257051
rect 20129 257023 20163 257051
rect 20191 257023 20239 257051
rect 19929 256989 20239 257023
rect 19929 256961 19977 256989
rect 20005 256961 20039 256989
rect 20067 256961 20101 256989
rect 20129 256961 20163 256989
rect 20191 256961 20239 256989
rect 19929 248175 20239 256961
rect 19929 248147 19977 248175
rect 20005 248147 20039 248175
rect 20067 248147 20101 248175
rect 20129 248147 20163 248175
rect 20191 248147 20239 248175
rect 19929 248113 20239 248147
rect 19929 248085 19977 248113
rect 20005 248085 20039 248113
rect 20067 248085 20101 248113
rect 20129 248085 20163 248113
rect 20191 248085 20239 248113
rect 19929 248051 20239 248085
rect 19929 248023 19977 248051
rect 20005 248023 20039 248051
rect 20067 248023 20101 248051
rect 20129 248023 20163 248051
rect 20191 248023 20239 248051
rect 19929 247989 20239 248023
rect 19929 247961 19977 247989
rect 20005 247961 20039 247989
rect 20067 247961 20101 247989
rect 20129 247961 20163 247989
rect 20191 247961 20239 247989
rect 19929 239175 20239 247961
rect 19929 239147 19977 239175
rect 20005 239147 20039 239175
rect 20067 239147 20101 239175
rect 20129 239147 20163 239175
rect 20191 239147 20239 239175
rect 19929 239113 20239 239147
rect 19929 239085 19977 239113
rect 20005 239085 20039 239113
rect 20067 239085 20101 239113
rect 20129 239085 20163 239113
rect 20191 239085 20239 239113
rect 19929 239051 20239 239085
rect 19929 239023 19977 239051
rect 20005 239023 20039 239051
rect 20067 239023 20101 239051
rect 20129 239023 20163 239051
rect 20191 239023 20239 239051
rect 19929 238989 20239 239023
rect 19929 238961 19977 238989
rect 20005 238961 20039 238989
rect 20067 238961 20101 238989
rect 20129 238961 20163 238989
rect 20191 238961 20239 238989
rect 19929 230175 20239 238961
rect 19929 230147 19977 230175
rect 20005 230147 20039 230175
rect 20067 230147 20101 230175
rect 20129 230147 20163 230175
rect 20191 230147 20239 230175
rect 19929 230113 20239 230147
rect 19929 230085 19977 230113
rect 20005 230085 20039 230113
rect 20067 230085 20101 230113
rect 20129 230085 20163 230113
rect 20191 230085 20239 230113
rect 19929 230051 20239 230085
rect 19929 230023 19977 230051
rect 20005 230023 20039 230051
rect 20067 230023 20101 230051
rect 20129 230023 20163 230051
rect 20191 230023 20239 230051
rect 19929 229989 20239 230023
rect 19929 229961 19977 229989
rect 20005 229961 20039 229989
rect 20067 229961 20101 229989
rect 20129 229961 20163 229989
rect 20191 229961 20239 229989
rect 19929 221175 20239 229961
rect 19929 221147 19977 221175
rect 20005 221147 20039 221175
rect 20067 221147 20101 221175
rect 20129 221147 20163 221175
rect 20191 221147 20239 221175
rect 19929 221113 20239 221147
rect 19929 221085 19977 221113
rect 20005 221085 20039 221113
rect 20067 221085 20101 221113
rect 20129 221085 20163 221113
rect 20191 221085 20239 221113
rect 19929 221051 20239 221085
rect 19929 221023 19977 221051
rect 20005 221023 20039 221051
rect 20067 221023 20101 221051
rect 20129 221023 20163 221051
rect 20191 221023 20239 221051
rect 19929 220989 20239 221023
rect 19929 220961 19977 220989
rect 20005 220961 20039 220989
rect 20067 220961 20101 220989
rect 20129 220961 20163 220989
rect 20191 220961 20239 220989
rect 19929 212175 20239 220961
rect 19929 212147 19977 212175
rect 20005 212147 20039 212175
rect 20067 212147 20101 212175
rect 20129 212147 20163 212175
rect 20191 212147 20239 212175
rect 19929 212113 20239 212147
rect 19929 212085 19977 212113
rect 20005 212085 20039 212113
rect 20067 212085 20101 212113
rect 20129 212085 20163 212113
rect 20191 212085 20239 212113
rect 19929 212051 20239 212085
rect 19929 212023 19977 212051
rect 20005 212023 20039 212051
rect 20067 212023 20101 212051
rect 20129 212023 20163 212051
rect 20191 212023 20239 212051
rect 19929 211989 20239 212023
rect 19929 211961 19977 211989
rect 20005 211961 20039 211989
rect 20067 211961 20101 211989
rect 20129 211961 20163 211989
rect 20191 211961 20239 211989
rect 19929 203175 20239 211961
rect 19929 203147 19977 203175
rect 20005 203147 20039 203175
rect 20067 203147 20101 203175
rect 20129 203147 20163 203175
rect 20191 203147 20239 203175
rect 19929 203113 20239 203147
rect 19929 203085 19977 203113
rect 20005 203085 20039 203113
rect 20067 203085 20101 203113
rect 20129 203085 20163 203113
rect 20191 203085 20239 203113
rect 19929 203051 20239 203085
rect 19929 203023 19977 203051
rect 20005 203023 20039 203051
rect 20067 203023 20101 203051
rect 20129 203023 20163 203051
rect 20191 203023 20239 203051
rect 19929 202989 20239 203023
rect 19929 202961 19977 202989
rect 20005 202961 20039 202989
rect 20067 202961 20101 202989
rect 20129 202961 20163 202989
rect 20191 202961 20239 202989
rect 19929 194175 20239 202961
rect 19929 194147 19977 194175
rect 20005 194147 20039 194175
rect 20067 194147 20101 194175
rect 20129 194147 20163 194175
rect 20191 194147 20239 194175
rect 19929 194113 20239 194147
rect 19929 194085 19977 194113
rect 20005 194085 20039 194113
rect 20067 194085 20101 194113
rect 20129 194085 20163 194113
rect 20191 194085 20239 194113
rect 19929 194051 20239 194085
rect 19929 194023 19977 194051
rect 20005 194023 20039 194051
rect 20067 194023 20101 194051
rect 20129 194023 20163 194051
rect 20191 194023 20239 194051
rect 19929 193989 20239 194023
rect 19929 193961 19977 193989
rect 20005 193961 20039 193989
rect 20067 193961 20101 193989
rect 20129 193961 20163 193989
rect 20191 193961 20239 193989
rect 19929 185175 20239 193961
rect 19929 185147 19977 185175
rect 20005 185147 20039 185175
rect 20067 185147 20101 185175
rect 20129 185147 20163 185175
rect 20191 185147 20239 185175
rect 19929 185113 20239 185147
rect 19929 185085 19977 185113
rect 20005 185085 20039 185113
rect 20067 185085 20101 185113
rect 20129 185085 20163 185113
rect 20191 185085 20239 185113
rect 19929 185051 20239 185085
rect 19929 185023 19977 185051
rect 20005 185023 20039 185051
rect 20067 185023 20101 185051
rect 20129 185023 20163 185051
rect 20191 185023 20239 185051
rect 19929 184989 20239 185023
rect 19929 184961 19977 184989
rect 20005 184961 20039 184989
rect 20067 184961 20101 184989
rect 20129 184961 20163 184989
rect 20191 184961 20239 184989
rect 19929 176175 20239 184961
rect 19929 176147 19977 176175
rect 20005 176147 20039 176175
rect 20067 176147 20101 176175
rect 20129 176147 20163 176175
rect 20191 176147 20239 176175
rect 19929 176113 20239 176147
rect 19929 176085 19977 176113
rect 20005 176085 20039 176113
rect 20067 176085 20101 176113
rect 20129 176085 20163 176113
rect 20191 176085 20239 176113
rect 19929 176051 20239 176085
rect 19929 176023 19977 176051
rect 20005 176023 20039 176051
rect 20067 176023 20101 176051
rect 20129 176023 20163 176051
rect 20191 176023 20239 176051
rect 19929 175989 20239 176023
rect 19929 175961 19977 175989
rect 20005 175961 20039 175989
rect 20067 175961 20101 175989
rect 20129 175961 20163 175989
rect 20191 175961 20239 175989
rect 19929 167175 20239 175961
rect 19929 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 20239 167175
rect 19929 167113 20239 167147
rect 19929 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 20239 167113
rect 19929 167051 20239 167085
rect 19929 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 20239 167051
rect 19929 166989 20239 167023
rect 19929 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 20239 166989
rect 19929 158175 20239 166961
rect 19929 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 20239 158175
rect 19929 158113 20239 158147
rect 19929 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 20239 158113
rect 19929 158051 20239 158085
rect 19929 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 20239 158051
rect 19929 157989 20239 158023
rect 19929 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 20239 157989
rect 19929 149175 20239 157961
rect 19929 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 20239 149175
rect 19929 149113 20239 149147
rect 19929 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 20239 149113
rect 19929 149051 20239 149085
rect 19929 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 20239 149051
rect 19929 148989 20239 149023
rect 19929 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 20239 148989
rect 19929 140175 20239 148961
rect 19929 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 20239 140175
rect 19929 140113 20239 140147
rect 19929 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 20239 140113
rect 19929 140051 20239 140085
rect 19929 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 20239 140051
rect 19929 139989 20239 140023
rect 19929 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 20239 139989
rect 19929 131175 20239 139961
rect 19929 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 20239 131175
rect 19929 131113 20239 131147
rect 19929 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 20239 131113
rect 19929 131051 20239 131085
rect 19929 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 20239 131051
rect 19929 130989 20239 131023
rect 19929 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 20239 130989
rect 19929 122175 20239 130961
rect 19929 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 20239 122175
rect 19929 122113 20239 122147
rect 19929 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 20239 122113
rect 19929 122051 20239 122085
rect 19929 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 20239 122051
rect 19929 121989 20239 122023
rect 19929 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 20239 121989
rect 19929 113175 20239 121961
rect 19929 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 20239 113175
rect 19929 113113 20239 113147
rect 19929 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 20239 113113
rect 19929 113051 20239 113085
rect 19929 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 20239 113051
rect 19929 112989 20239 113023
rect 19929 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 20239 112989
rect 19929 104175 20239 112961
rect 19929 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 20239 104175
rect 19929 104113 20239 104147
rect 19929 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 20239 104113
rect 19929 104051 20239 104085
rect 19929 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 20239 104051
rect 19929 103989 20239 104023
rect 19929 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 20239 103989
rect 19929 95175 20239 103961
rect 19929 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 20239 95175
rect 19929 95113 20239 95147
rect 19929 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 20239 95113
rect 19929 95051 20239 95085
rect 19929 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 20239 95051
rect 19929 94989 20239 95023
rect 19929 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 20239 94989
rect 19929 86175 20239 94961
rect 19929 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 20239 86175
rect 19929 86113 20239 86147
rect 19929 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 20239 86113
rect 19929 86051 20239 86085
rect 19929 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 20239 86051
rect 19929 85989 20239 86023
rect 19929 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 20239 85989
rect 19929 77175 20239 85961
rect 19929 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 20239 77175
rect 19929 77113 20239 77147
rect 19929 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 20239 77113
rect 19929 77051 20239 77085
rect 19929 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 20239 77051
rect 19929 76989 20239 77023
rect 19929 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 20239 76989
rect 19929 68175 20239 76961
rect 19929 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 20239 68175
rect 19929 68113 20239 68147
rect 19929 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 20239 68113
rect 19929 68051 20239 68085
rect 19929 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 20239 68051
rect 19929 67989 20239 68023
rect 19929 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 20239 67989
rect 19929 59175 20239 67961
rect 19929 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 20239 59175
rect 19929 59113 20239 59147
rect 19929 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 20239 59113
rect 19929 59051 20239 59085
rect 19929 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 20239 59051
rect 19929 58989 20239 59023
rect 19929 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 20239 58989
rect 19929 50175 20239 58961
rect 19929 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 20239 50175
rect 19929 50113 20239 50147
rect 19929 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 20239 50113
rect 19929 50051 20239 50085
rect 19929 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 20239 50051
rect 19929 49989 20239 50023
rect 19929 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 20239 49989
rect 19929 41175 20239 49961
rect 19929 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 20239 41175
rect 19929 41113 20239 41147
rect 19929 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 20239 41113
rect 19929 41051 20239 41085
rect 19929 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 20239 41051
rect 19929 40989 20239 41023
rect 19929 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 20239 40989
rect 19929 32175 20239 40961
rect 19929 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 20239 32175
rect 19929 32113 20239 32147
rect 19929 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 20239 32113
rect 19929 32051 20239 32085
rect 19929 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 20239 32051
rect 19929 31989 20239 32023
rect 19929 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 20239 31989
rect 19929 23175 20239 31961
rect 19929 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 20239 23175
rect 19929 23113 20239 23147
rect 19929 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 20239 23113
rect 19929 23051 20239 23085
rect 19929 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 20239 23051
rect 19929 22989 20239 23023
rect 19929 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 20239 22989
rect 19929 14175 20239 22961
rect 19929 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 20239 14175
rect 19929 14113 20239 14147
rect 19929 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 20239 14113
rect 19929 14051 20239 14085
rect 19929 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 20239 14051
rect 19929 13989 20239 14023
rect 19929 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 20239 13989
rect 19929 5175 20239 13961
rect 19929 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 20239 5175
rect 19929 5113 20239 5147
rect 19929 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 20239 5113
rect 19929 5051 20239 5085
rect 19929 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 20239 5051
rect 19929 4989 20239 5023
rect 19929 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 20239 4989
rect 19929 -560 20239 4961
rect 19929 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 20239 -560
rect 19929 -622 20239 -588
rect 19929 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 20239 -622
rect 19929 -684 20239 -650
rect 19929 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 20239 -684
rect 19929 -746 20239 -712
rect 19929 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 20239 -746
rect 19929 -822 20239 -774
rect 33429 298606 33739 299134
rect 33429 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 33739 298606
rect 33429 298544 33739 298578
rect 33429 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 33739 298544
rect 33429 298482 33739 298516
rect 33429 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 33739 298482
rect 33429 298420 33739 298454
rect 33429 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 33739 298420
rect 33429 290175 33739 298392
rect 33429 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 33739 290175
rect 33429 290113 33739 290147
rect 33429 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 33739 290113
rect 33429 290051 33739 290085
rect 33429 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 33739 290051
rect 33429 289989 33739 290023
rect 33429 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 33739 289989
rect 33429 281175 33739 289961
rect 33429 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 33739 281175
rect 33429 281113 33739 281147
rect 33429 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 33739 281113
rect 33429 281051 33739 281085
rect 33429 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 33739 281051
rect 33429 280989 33739 281023
rect 33429 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 33739 280989
rect 33429 272175 33739 280961
rect 33429 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 33739 272175
rect 33429 272113 33739 272147
rect 33429 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 33739 272113
rect 33429 272051 33739 272085
rect 33429 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 33739 272051
rect 33429 271989 33739 272023
rect 33429 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 33739 271989
rect 33429 263175 33739 271961
rect 33429 263147 33477 263175
rect 33505 263147 33539 263175
rect 33567 263147 33601 263175
rect 33629 263147 33663 263175
rect 33691 263147 33739 263175
rect 33429 263113 33739 263147
rect 33429 263085 33477 263113
rect 33505 263085 33539 263113
rect 33567 263085 33601 263113
rect 33629 263085 33663 263113
rect 33691 263085 33739 263113
rect 33429 263051 33739 263085
rect 33429 263023 33477 263051
rect 33505 263023 33539 263051
rect 33567 263023 33601 263051
rect 33629 263023 33663 263051
rect 33691 263023 33739 263051
rect 33429 262989 33739 263023
rect 33429 262961 33477 262989
rect 33505 262961 33539 262989
rect 33567 262961 33601 262989
rect 33629 262961 33663 262989
rect 33691 262961 33739 262989
rect 33429 254175 33739 262961
rect 33429 254147 33477 254175
rect 33505 254147 33539 254175
rect 33567 254147 33601 254175
rect 33629 254147 33663 254175
rect 33691 254147 33739 254175
rect 33429 254113 33739 254147
rect 33429 254085 33477 254113
rect 33505 254085 33539 254113
rect 33567 254085 33601 254113
rect 33629 254085 33663 254113
rect 33691 254085 33739 254113
rect 33429 254051 33739 254085
rect 33429 254023 33477 254051
rect 33505 254023 33539 254051
rect 33567 254023 33601 254051
rect 33629 254023 33663 254051
rect 33691 254023 33739 254051
rect 33429 253989 33739 254023
rect 33429 253961 33477 253989
rect 33505 253961 33539 253989
rect 33567 253961 33601 253989
rect 33629 253961 33663 253989
rect 33691 253961 33739 253989
rect 33429 245175 33739 253961
rect 33429 245147 33477 245175
rect 33505 245147 33539 245175
rect 33567 245147 33601 245175
rect 33629 245147 33663 245175
rect 33691 245147 33739 245175
rect 33429 245113 33739 245147
rect 33429 245085 33477 245113
rect 33505 245085 33539 245113
rect 33567 245085 33601 245113
rect 33629 245085 33663 245113
rect 33691 245085 33739 245113
rect 33429 245051 33739 245085
rect 33429 245023 33477 245051
rect 33505 245023 33539 245051
rect 33567 245023 33601 245051
rect 33629 245023 33663 245051
rect 33691 245023 33739 245051
rect 33429 244989 33739 245023
rect 33429 244961 33477 244989
rect 33505 244961 33539 244989
rect 33567 244961 33601 244989
rect 33629 244961 33663 244989
rect 33691 244961 33739 244989
rect 33429 236175 33739 244961
rect 33429 236147 33477 236175
rect 33505 236147 33539 236175
rect 33567 236147 33601 236175
rect 33629 236147 33663 236175
rect 33691 236147 33739 236175
rect 33429 236113 33739 236147
rect 33429 236085 33477 236113
rect 33505 236085 33539 236113
rect 33567 236085 33601 236113
rect 33629 236085 33663 236113
rect 33691 236085 33739 236113
rect 33429 236051 33739 236085
rect 33429 236023 33477 236051
rect 33505 236023 33539 236051
rect 33567 236023 33601 236051
rect 33629 236023 33663 236051
rect 33691 236023 33739 236051
rect 33429 235989 33739 236023
rect 33429 235961 33477 235989
rect 33505 235961 33539 235989
rect 33567 235961 33601 235989
rect 33629 235961 33663 235989
rect 33691 235961 33739 235989
rect 33429 227175 33739 235961
rect 33429 227147 33477 227175
rect 33505 227147 33539 227175
rect 33567 227147 33601 227175
rect 33629 227147 33663 227175
rect 33691 227147 33739 227175
rect 33429 227113 33739 227147
rect 33429 227085 33477 227113
rect 33505 227085 33539 227113
rect 33567 227085 33601 227113
rect 33629 227085 33663 227113
rect 33691 227085 33739 227113
rect 33429 227051 33739 227085
rect 33429 227023 33477 227051
rect 33505 227023 33539 227051
rect 33567 227023 33601 227051
rect 33629 227023 33663 227051
rect 33691 227023 33739 227051
rect 33429 226989 33739 227023
rect 33429 226961 33477 226989
rect 33505 226961 33539 226989
rect 33567 226961 33601 226989
rect 33629 226961 33663 226989
rect 33691 226961 33739 226989
rect 33429 218175 33739 226961
rect 33429 218147 33477 218175
rect 33505 218147 33539 218175
rect 33567 218147 33601 218175
rect 33629 218147 33663 218175
rect 33691 218147 33739 218175
rect 33429 218113 33739 218147
rect 33429 218085 33477 218113
rect 33505 218085 33539 218113
rect 33567 218085 33601 218113
rect 33629 218085 33663 218113
rect 33691 218085 33739 218113
rect 33429 218051 33739 218085
rect 33429 218023 33477 218051
rect 33505 218023 33539 218051
rect 33567 218023 33601 218051
rect 33629 218023 33663 218051
rect 33691 218023 33739 218051
rect 33429 217989 33739 218023
rect 33429 217961 33477 217989
rect 33505 217961 33539 217989
rect 33567 217961 33601 217989
rect 33629 217961 33663 217989
rect 33691 217961 33739 217989
rect 33429 209175 33739 217961
rect 33429 209147 33477 209175
rect 33505 209147 33539 209175
rect 33567 209147 33601 209175
rect 33629 209147 33663 209175
rect 33691 209147 33739 209175
rect 33429 209113 33739 209147
rect 33429 209085 33477 209113
rect 33505 209085 33539 209113
rect 33567 209085 33601 209113
rect 33629 209085 33663 209113
rect 33691 209085 33739 209113
rect 33429 209051 33739 209085
rect 33429 209023 33477 209051
rect 33505 209023 33539 209051
rect 33567 209023 33601 209051
rect 33629 209023 33663 209051
rect 33691 209023 33739 209051
rect 33429 208989 33739 209023
rect 33429 208961 33477 208989
rect 33505 208961 33539 208989
rect 33567 208961 33601 208989
rect 33629 208961 33663 208989
rect 33691 208961 33739 208989
rect 33429 200175 33739 208961
rect 33429 200147 33477 200175
rect 33505 200147 33539 200175
rect 33567 200147 33601 200175
rect 33629 200147 33663 200175
rect 33691 200147 33739 200175
rect 33429 200113 33739 200147
rect 33429 200085 33477 200113
rect 33505 200085 33539 200113
rect 33567 200085 33601 200113
rect 33629 200085 33663 200113
rect 33691 200085 33739 200113
rect 33429 200051 33739 200085
rect 33429 200023 33477 200051
rect 33505 200023 33539 200051
rect 33567 200023 33601 200051
rect 33629 200023 33663 200051
rect 33691 200023 33739 200051
rect 33429 199989 33739 200023
rect 33429 199961 33477 199989
rect 33505 199961 33539 199989
rect 33567 199961 33601 199989
rect 33629 199961 33663 199989
rect 33691 199961 33739 199989
rect 33429 191175 33739 199961
rect 33429 191147 33477 191175
rect 33505 191147 33539 191175
rect 33567 191147 33601 191175
rect 33629 191147 33663 191175
rect 33691 191147 33739 191175
rect 33429 191113 33739 191147
rect 33429 191085 33477 191113
rect 33505 191085 33539 191113
rect 33567 191085 33601 191113
rect 33629 191085 33663 191113
rect 33691 191085 33739 191113
rect 33429 191051 33739 191085
rect 33429 191023 33477 191051
rect 33505 191023 33539 191051
rect 33567 191023 33601 191051
rect 33629 191023 33663 191051
rect 33691 191023 33739 191051
rect 33429 190989 33739 191023
rect 33429 190961 33477 190989
rect 33505 190961 33539 190989
rect 33567 190961 33601 190989
rect 33629 190961 33663 190989
rect 33691 190961 33739 190989
rect 33429 182175 33739 190961
rect 33429 182147 33477 182175
rect 33505 182147 33539 182175
rect 33567 182147 33601 182175
rect 33629 182147 33663 182175
rect 33691 182147 33739 182175
rect 33429 182113 33739 182147
rect 33429 182085 33477 182113
rect 33505 182085 33539 182113
rect 33567 182085 33601 182113
rect 33629 182085 33663 182113
rect 33691 182085 33739 182113
rect 33429 182051 33739 182085
rect 33429 182023 33477 182051
rect 33505 182023 33539 182051
rect 33567 182023 33601 182051
rect 33629 182023 33663 182051
rect 33691 182023 33739 182051
rect 33429 181989 33739 182023
rect 33429 181961 33477 181989
rect 33505 181961 33539 181989
rect 33567 181961 33601 181989
rect 33629 181961 33663 181989
rect 33691 181961 33739 181989
rect 33429 173175 33739 181961
rect 33429 173147 33477 173175
rect 33505 173147 33539 173175
rect 33567 173147 33601 173175
rect 33629 173147 33663 173175
rect 33691 173147 33739 173175
rect 33429 173113 33739 173147
rect 33429 173085 33477 173113
rect 33505 173085 33539 173113
rect 33567 173085 33601 173113
rect 33629 173085 33663 173113
rect 33691 173085 33739 173113
rect 33429 173051 33739 173085
rect 33429 173023 33477 173051
rect 33505 173023 33539 173051
rect 33567 173023 33601 173051
rect 33629 173023 33663 173051
rect 33691 173023 33739 173051
rect 33429 172989 33739 173023
rect 33429 172961 33477 172989
rect 33505 172961 33539 172989
rect 33567 172961 33601 172989
rect 33629 172961 33663 172989
rect 33691 172961 33739 172989
rect 33429 164175 33739 172961
rect 33429 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 33739 164175
rect 33429 164113 33739 164147
rect 33429 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 33739 164113
rect 33429 164051 33739 164085
rect 33429 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 33739 164051
rect 33429 163989 33739 164023
rect 33429 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 33739 163989
rect 33429 155175 33739 163961
rect 33429 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 33739 155175
rect 33429 155113 33739 155147
rect 33429 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 33739 155113
rect 33429 155051 33739 155085
rect 33429 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 33739 155051
rect 33429 154989 33739 155023
rect 33429 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 33739 154989
rect 33429 146175 33739 154961
rect 33429 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 33739 146175
rect 33429 146113 33739 146147
rect 33429 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 33739 146113
rect 33429 146051 33739 146085
rect 33429 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 33739 146051
rect 33429 145989 33739 146023
rect 33429 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 33739 145989
rect 33429 137175 33739 145961
rect 33429 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 33739 137175
rect 33429 137113 33739 137147
rect 33429 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 33739 137113
rect 33429 137051 33739 137085
rect 33429 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 33739 137051
rect 33429 136989 33739 137023
rect 33429 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 33739 136989
rect 33429 128175 33739 136961
rect 33429 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 33739 128175
rect 33429 128113 33739 128147
rect 33429 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 33739 128113
rect 33429 128051 33739 128085
rect 33429 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 33739 128051
rect 33429 127989 33739 128023
rect 33429 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 33739 127989
rect 33429 119175 33739 127961
rect 33429 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 33739 119175
rect 33429 119113 33739 119147
rect 33429 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 33739 119113
rect 33429 119051 33739 119085
rect 33429 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 33739 119051
rect 33429 118989 33739 119023
rect 33429 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 33739 118989
rect 33429 110175 33739 118961
rect 33429 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 33739 110175
rect 33429 110113 33739 110147
rect 33429 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 33739 110113
rect 33429 110051 33739 110085
rect 33429 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 33739 110051
rect 33429 109989 33739 110023
rect 33429 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 33739 109989
rect 33429 101175 33739 109961
rect 33429 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 33739 101175
rect 33429 101113 33739 101147
rect 33429 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 33739 101113
rect 33429 101051 33739 101085
rect 33429 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 33739 101051
rect 33429 100989 33739 101023
rect 33429 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 33739 100989
rect 33429 92175 33739 100961
rect 33429 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 33739 92175
rect 33429 92113 33739 92147
rect 33429 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 33739 92113
rect 33429 92051 33739 92085
rect 33429 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 33739 92051
rect 33429 91989 33739 92023
rect 33429 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 33739 91989
rect 33429 83175 33739 91961
rect 33429 83147 33477 83175
rect 33505 83147 33539 83175
rect 33567 83147 33601 83175
rect 33629 83147 33663 83175
rect 33691 83147 33739 83175
rect 33429 83113 33739 83147
rect 33429 83085 33477 83113
rect 33505 83085 33539 83113
rect 33567 83085 33601 83113
rect 33629 83085 33663 83113
rect 33691 83085 33739 83113
rect 33429 83051 33739 83085
rect 33429 83023 33477 83051
rect 33505 83023 33539 83051
rect 33567 83023 33601 83051
rect 33629 83023 33663 83051
rect 33691 83023 33739 83051
rect 33429 82989 33739 83023
rect 33429 82961 33477 82989
rect 33505 82961 33539 82989
rect 33567 82961 33601 82989
rect 33629 82961 33663 82989
rect 33691 82961 33739 82989
rect 33429 74175 33739 82961
rect 33429 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 33739 74175
rect 33429 74113 33739 74147
rect 33429 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 33739 74113
rect 33429 74051 33739 74085
rect 33429 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 33739 74051
rect 33429 73989 33739 74023
rect 33429 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 33739 73989
rect 33429 65175 33739 73961
rect 33429 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 33739 65175
rect 33429 65113 33739 65147
rect 33429 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 33739 65113
rect 33429 65051 33739 65085
rect 33429 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 33739 65051
rect 33429 64989 33739 65023
rect 33429 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 33739 64989
rect 33429 56175 33739 64961
rect 33429 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 33739 56175
rect 33429 56113 33739 56147
rect 33429 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 33739 56113
rect 33429 56051 33739 56085
rect 33429 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 33739 56051
rect 33429 55989 33739 56023
rect 33429 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 33739 55989
rect 33429 47175 33739 55961
rect 33429 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 33739 47175
rect 33429 47113 33739 47147
rect 33429 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 33739 47113
rect 33429 47051 33739 47085
rect 33429 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 33739 47051
rect 33429 46989 33739 47023
rect 33429 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 33739 46989
rect 33429 38175 33739 46961
rect 33429 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 33739 38175
rect 33429 38113 33739 38147
rect 33429 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 33739 38113
rect 33429 38051 33739 38085
rect 33429 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 33739 38051
rect 33429 37989 33739 38023
rect 33429 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 33739 37989
rect 33429 29175 33739 37961
rect 33429 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 33739 29175
rect 33429 29113 33739 29147
rect 33429 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 33739 29113
rect 33429 29051 33739 29085
rect 33429 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 33739 29051
rect 33429 28989 33739 29023
rect 33429 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 33739 28989
rect 33429 20175 33739 28961
rect 33429 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 33739 20175
rect 33429 20113 33739 20147
rect 33429 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 33739 20113
rect 33429 20051 33739 20085
rect 33429 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 33739 20051
rect 33429 19989 33739 20023
rect 33429 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 33739 19989
rect 33429 11175 33739 19961
rect 33429 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 33739 11175
rect 33429 11113 33739 11147
rect 33429 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 33739 11113
rect 33429 11051 33739 11085
rect 33429 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 33739 11051
rect 33429 10989 33739 11023
rect 33429 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 33739 10989
rect 33429 2175 33739 10961
rect 33429 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 33739 2175
rect 33429 2113 33739 2147
rect 33429 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 33739 2113
rect 33429 2051 33739 2085
rect 33429 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 33739 2051
rect 33429 1989 33739 2023
rect 33429 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 33739 1989
rect 33429 -80 33739 1961
rect 33429 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 33739 -80
rect 33429 -142 33739 -108
rect 33429 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 33739 -142
rect 33429 -204 33739 -170
rect 33429 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 33739 -204
rect 33429 -266 33739 -232
rect 33429 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 33739 -266
rect 33429 -822 33739 -294
rect 35289 299086 35599 299134
rect 35289 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 35599 299086
rect 35289 299024 35599 299058
rect 35289 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 35599 299024
rect 35289 298962 35599 298996
rect 35289 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 35599 298962
rect 35289 298900 35599 298934
rect 35289 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 35599 298900
rect 35289 293175 35599 298872
rect 35289 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 35599 293175
rect 35289 293113 35599 293147
rect 35289 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 35599 293113
rect 35289 293051 35599 293085
rect 35289 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 35599 293051
rect 35289 292989 35599 293023
rect 35289 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 35599 292989
rect 35289 284175 35599 292961
rect 35289 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 35599 284175
rect 35289 284113 35599 284147
rect 35289 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 35599 284113
rect 35289 284051 35599 284085
rect 35289 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 35599 284051
rect 35289 283989 35599 284023
rect 35289 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 35599 283989
rect 35289 275175 35599 283961
rect 35289 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 35599 275175
rect 35289 275113 35599 275147
rect 35289 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 35599 275113
rect 35289 275051 35599 275085
rect 35289 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 35599 275051
rect 35289 274989 35599 275023
rect 35289 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 35599 274989
rect 35289 266175 35599 274961
rect 35289 266147 35337 266175
rect 35365 266147 35399 266175
rect 35427 266147 35461 266175
rect 35489 266147 35523 266175
rect 35551 266147 35599 266175
rect 35289 266113 35599 266147
rect 35289 266085 35337 266113
rect 35365 266085 35399 266113
rect 35427 266085 35461 266113
rect 35489 266085 35523 266113
rect 35551 266085 35599 266113
rect 35289 266051 35599 266085
rect 35289 266023 35337 266051
rect 35365 266023 35399 266051
rect 35427 266023 35461 266051
rect 35489 266023 35523 266051
rect 35551 266023 35599 266051
rect 35289 265989 35599 266023
rect 35289 265961 35337 265989
rect 35365 265961 35399 265989
rect 35427 265961 35461 265989
rect 35489 265961 35523 265989
rect 35551 265961 35599 265989
rect 35289 257175 35599 265961
rect 35289 257147 35337 257175
rect 35365 257147 35399 257175
rect 35427 257147 35461 257175
rect 35489 257147 35523 257175
rect 35551 257147 35599 257175
rect 35289 257113 35599 257147
rect 35289 257085 35337 257113
rect 35365 257085 35399 257113
rect 35427 257085 35461 257113
rect 35489 257085 35523 257113
rect 35551 257085 35599 257113
rect 35289 257051 35599 257085
rect 35289 257023 35337 257051
rect 35365 257023 35399 257051
rect 35427 257023 35461 257051
rect 35489 257023 35523 257051
rect 35551 257023 35599 257051
rect 35289 256989 35599 257023
rect 35289 256961 35337 256989
rect 35365 256961 35399 256989
rect 35427 256961 35461 256989
rect 35489 256961 35523 256989
rect 35551 256961 35599 256989
rect 35289 248175 35599 256961
rect 35289 248147 35337 248175
rect 35365 248147 35399 248175
rect 35427 248147 35461 248175
rect 35489 248147 35523 248175
rect 35551 248147 35599 248175
rect 35289 248113 35599 248147
rect 35289 248085 35337 248113
rect 35365 248085 35399 248113
rect 35427 248085 35461 248113
rect 35489 248085 35523 248113
rect 35551 248085 35599 248113
rect 35289 248051 35599 248085
rect 35289 248023 35337 248051
rect 35365 248023 35399 248051
rect 35427 248023 35461 248051
rect 35489 248023 35523 248051
rect 35551 248023 35599 248051
rect 35289 247989 35599 248023
rect 35289 247961 35337 247989
rect 35365 247961 35399 247989
rect 35427 247961 35461 247989
rect 35489 247961 35523 247989
rect 35551 247961 35599 247989
rect 35289 239175 35599 247961
rect 35289 239147 35337 239175
rect 35365 239147 35399 239175
rect 35427 239147 35461 239175
rect 35489 239147 35523 239175
rect 35551 239147 35599 239175
rect 35289 239113 35599 239147
rect 35289 239085 35337 239113
rect 35365 239085 35399 239113
rect 35427 239085 35461 239113
rect 35489 239085 35523 239113
rect 35551 239085 35599 239113
rect 35289 239051 35599 239085
rect 35289 239023 35337 239051
rect 35365 239023 35399 239051
rect 35427 239023 35461 239051
rect 35489 239023 35523 239051
rect 35551 239023 35599 239051
rect 35289 238989 35599 239023
rect 35289 238961 35337 238989
rect 35365 238961 35399 238989
rect 35427 238961 35461 238989
rect 35489 238961 35523 238989
rect 35551 238961 35599 238989
rect 35289 230175 35599 238961
rect 35289 230147 35337 230175
rect 35365 230147 35399 230175
rect 35427 230147 35461 230175
rect 35489 230147 35523 230175
rect 35551 230147 35599 230175
rect 35289 230113 35599 230147
rect 35289 230085 35337 230113
rect 35365 230085 35399 230113
rect 35427 230085 35461 230113
rect 35489 230085 35523 230113
rect 35551 230085 35599 230113
rect 35289 230051 35599 230085
rect 35289 230023 35337 230051
rect 35365 230023 35399 230051
rect 35427 230023 35461 230051
rect 35489 230023 35523 230051
rect 35551 230023 35599 230051
rect 35289 229989 35599 230023
rect 35289 229961 35337 229989
rect 35365 229961 35399 229989
rect 35427 229961 35461 229989
rect 35489 229961 35523 229989
rect 35551 229961 35599 229989
rect 35289 221175 35599 229961
rect 35289 221147 35337 221175
rect 35365 221147 35399 221175
rect 35427 221147 35461 221175
rect 35489 221147 35523 221175
rect 35551 221147 35599 221175
rect 35289 221113 35599 221147
rect 35289 221085 35337 221113
rect 35365 221085 35399 221113
rect 35427 221085 35461 221113
rect 35489 221085 35523 221113
rect 35551 221085 35599 221113
rect 35289 221051 35599 221085
rect 35289 221023 35337 221051
rect 35365 221023 35399 221051
rect 35427 221023 35461 221051
rect 35489 221023 35523 221051
rect 35551 221023 35599 221051
rect 35289 220989 35599 221023
rect 35289 220961 35337 220989
rect 35365 220961 35399 220989
rect 35427 220961 35461 220989
rect 35489 220961 35523 220989
rect 35551 220961 35599 220989
rect 35289 212175 35599 220961
rect 35289 212147 35337 212175
rect 35365 212147 35399 212175
rect 35427 212147 35461 212175
rect 35489 212147 35523 212175
rect 35551 212147 35599 212175
rect 35289 212113 35599 212147
rect 35289 212085 35337 212113
rect 35365 212085 35399 212113
rect 35427 212085 35461 212113
rect 35489 212085 35523 212113
rect 35551 212085 35599 212113
rect 35289 212051 35599 212085
rect 35289 212023 35337 212051
rect 35365 212023 35399 212051
rect 35427 212023 35461 212051
rect 35489 212023 35523 212051
rect 35551 212023 35599 212051
rect 35289 211989 35599 212023
rect 35289 211961 35337 211989
rect 35365 211961 35399 211989
rect 35427 211961 35461 211989
rect 35489 211961 35523 211989
rect 35551 211961 35599 211989
rect 35289 203175 35599 211961
rect 35289 203147 35337 203175
rect 35365 203147 35399 203175
rect 35427 203147 35461 203175
rect 35489 203147 35523 203175
rect 35551 203147 35599 203175
rect 35289 203113 35599 203147
rect 35289 203085 35337 203113
rect 35365 203085 35399 203113
rect 35427 203085 35461 203113
rect 35489 203085 35523 203113
rect 35551 203085 35599 203113
rect 35289 203051 35599 203085
rect 35289 203023 35337 203051
rect 35365 203023 35399 203051
rect 35427 203023 35461 203051
rect 35489 203023 35523 203051
rect 35551 203023 35599 203051
rect 35289 202989 35599 203023
rect 35289 202961 35337 202989
rect 35365 202961 35399 202989
rect 35427 202961 35461 202989
rect 35489 202961 35523 202989
rect 35551 202961 35599 202989
rect 35289 194175 35599 202961
rect 35289 194147 35337 194175
rect 35365 194147 35399 194175
rect 35427 194147 35461 194175
rect 35489 194147 35523 194175
rect 35551 194147 35599 194175
rect 35289 194113 35599 194147
rect 35289 194085 35337 194113
rect 35365 194085 35399 194113
rect 35427 194085 35461 194113
rect 35489 194085 35523 194113
rect 35551 194085 35599 194113
rect 35289 194051 35599 194085
rect 35289 194023 35337 194051
rect 35365 194023 35399 194051
rect 35427 194023 35461 194051
rect 35489 194023 35523 194051
rect 35551 194023 35599 194051
rect 35289 193989 35599 194023
rect 35289 193961 35337 193989
rect 35365 193961 35399 193989
rect 35427 193961 35461 193989
rect 35489 193961 35523 193989
rect 35551 193961 35599 193989
rect 35289 185175 35599 193961
rect 35289 185147 35337 185175
rect 35365 185147 35399 185175
rect 35427 185147 35461 185175
rect 35489 185147 35523 185175
rect 35551 185147 35599 185175
rect 35289 185113 35599 185147
rect 35289 185085 35337 185113
rect 35365 185085 35399 185113
rect 35427 185085 35461 185113
rect 35489 185085 35523 185113
rect 35551 185085 35599 185113
rect 35289 185051 35599 185085
rect 35289 185023 35337 185051
rect 35365 185023 35399 185051
rect 35427 185023 35461 185051
rect 35489 185023 35523 185051
rect 35551 185023 35599 185051
rect 35289 184989 35599 185023
rect 35289 184961 35337 184989
rect 35365 184961 35399 184989
rect 35427 184961 35461 184989
rect 35489 184961 35523 184989
rect 35551 184961 35599 184989
rect 35289 176175 35599 184961
rect 35289 176147 35337 176175
rect 35365 176147 35399 176175
rect 35427 176147 35461 176175
rect 35489 176147 35523 176175
rect 35551 176147 35599 176175
rect 35289 176113 35599 176147
rect 35289 176085 35337 176113
rect 35365 176085 35399 176113
rect 35427 176085 35461 176113
rect 35489 176085 35523 176113
rect 35551 176085 35599 176113
rect 35289 176051 35599 176085
rect 35289 176023 35337 176051
rect 35365 176023 35399 176051
rect 35427 176023 35461 176051
rect 35489 176023 35523 176051
rect 35551 176023 35599 176051
rect 35289 175989 35599 176023
rect 35289 175961 35337 175989
rect 35365 175961 35399 175989
rect 35427 175961 35461 175989
rect 35489 175961 35523 175989
rect 35551 175961 35599 175989
rect 35289 167175 35599 175961
rect 35289 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 35599 167175
rect 35289 167113 35599 167147
rect 35289 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 35599 167113
rect 35289 167051 35599 167085
rect 35289 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 35599 167051
rect 35289 166989 35599 167023
rect 35289 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 35599 166989
rect 35289 158175 35599 166961
rect 35289 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 35599 158175
rect 35289 158113 35599 158147
rect 35289 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 35599 158113
rect 35289 158051 35599 158085
rect 35289 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 35599 158051
rect 35289 157989 35599 158023
rect 35289 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 35599 157989
rect 35289 149175 35599 157961
rect 35289 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 35599 149175
rect 35289 149113 35599 149147
rect 35289 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 35599 149113
rect 35289 149051 35599 149085
rect 35289 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 35599 149051
rect 35289 148989 35599 149023
rect 35289 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 35599 148989
rect 35289 140175 35599 148961
rect 35289 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 35599 140175
rect 35289 140113 35599 140147
rect 35289 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 35599 140113
rect 35289 140051 35599 140085
rect 35289 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 35599 140051
rect 35289 139989 35599 140023
rect 35289 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 35599 139989
rect 35289 131175 35599 139961
rect 35289 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 35599 131175
rect 35289 131113 35599 131147
rect 35289 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 35599 131113
rect 35289 131051 35599 131085
rect 35289 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 35599 131051
rect 35289 130989 35599 131023
rect 35289 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 35599 130989
rect 35289 122175 35599 130961
rect 35289 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 35599 122175
rect 35289 122113 35599 122147
rect 35289 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 35599 122113
rect 35289 122051 35599 122085
rect 35289 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 35599 122051
rect 35289 121989 35599 122023
rect 35289 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 35599 121989
rect 35289 113175 35599 121961
rect 35289 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 35599 113175
rect 35289 113113 35599 113147
rect 35289 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 35599 113113
rect 35289 113051 35599 113085
rect 35289 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 35599 113051
rect 35289 112989 35599 113023
rect 35289 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 35599 112989
rect 35289 104175 35599 112961
rect 35289 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 35599 104175
rect 35289 104113 35599 104147
rect 35289 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 35599 104113
rect 35289 104051 35599 104085
rect 35289 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 35599 104051
rect 35289 103989 35599 104023
rect 35289 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 35599 103989
rect 35289 95175 35599 103961
rect 35289 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 35599 95175
rect 35289 95113 35599 95147
rect 35289 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 35599 95113
rect 35289 95051 35599 95085
rect 35289 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 35599 95051
rect 35289 94989 35599 95023
rect 35289 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 35599 94989
rect 35289 86175 35599 94961
rect 35289 86147 35337 86175
rect 35365 86147 35399 86175
rect 35427 86147 35461 86175
rect 35489 86147 35523 86175
rect 35551 86147 35599 86175
rect 35289 86113 35599 86147
rect 35289 86085 35337 86113
rect 35365 86085 35399 86113
rect 35427 86085 35461 86113
rect 35489 86085 35523 86113
rect 35551 86085 35599 86113
rect 35289 86051 35599 86085
rect 35289 86023 35337 86051
rect 35365 86023 35399 86051
rect 35427 86023 35461 86051
rect 35489 86023 35523 86051
rect 35551 86023 35599 86051
rect 35289 85989 35599 86023
rect 35289 85961 35337 85989
rect 35365 85961 35399 85989
rect 35427 85961 35461 85989
rect 35489 85961 35523 85989
rect 35551 85961 35599 85989
rect 35289 77175 35599 85961
rect 35289 77147 35337 77175
rect 35365 77147 35399 77175
rect 35427 77147 35461 77175
rect 35489 77147 35523 77175
rect 35551 77147 35599 77175
rect 35289 77113 35599 77147
rect 35289 77085 35337 77113
rect 35365 77085 35399 77113
rect 35427 77085 35461 77113
rect 35489 77085 35523 77113
rect 35551 77085 35599 77113
rect 35289 77051 35599 77085
rect 35289 77023 35337 77051
rect 35365 77023 35399 77051
rect 35427 77023 35461 77051
rect 35489 77023 35523 77051
rect 35551 77023 35599 77051
rect 35289 76989 35599 77023
rect 35289 76961 35337 76989
rect 35365 76961 35399 76989
rect 35427 76961 35461 76989
rect 35489 76961 35523 76989
rect 35551 76961 35599 76989
rect 35289 68175 35599 76961
rect 35289 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 35599 68175
rect 35289 68113 35599 68147
rect 35289 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 35599 68113
rect 35289 68051 35599 68085
rect 35289 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 35599 68051
rect 35289 67989 35599 68023
rect 35289 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 35599 67989
rect 35289 59175 35599 67961
rect 35289 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 35599 59175
rect 35289 59113 35599 59147
rect 35289 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 35599 59113
rect 35289 59051 35599 59085
rect 35289 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 35599 59051
rect 35289 58989 35599 59023
rect 35289 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 35599 58989
rect 35289 50175 35599 58961
rect 35289 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 35599 50175
rect 35289 50113 35599 50147
rect 35289 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 35599 50113
rect 35289 50051 35599 50085
rect 35289 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 35599 50051
rect 35289 49989 35599 50023
rect 35289 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 35599 49989
rect 35289 41175 35599 49961
rect 35289 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 35599 41175
rect 35289 41113 35599 41147
rect 35289 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 35599 41113
rect 35289 41051 35599 41085
rect 35289 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 35599 41051
rect 35289 40989 35599 41023
rect 35289 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 35599 40989
rect 35289 32175 35599 40961
rect 35289 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 35599 32175
rect 35289 32113 35599 32147
rect 35289 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 35599 32113
rect 35289 32051 35599 32085
rect 35289 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 35599 32051
rect 35289 31989 35599 32023
rect 35289 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 35599 31989
rect 35289 23175 35599 31961
rect 35289 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 35599 23175
rect 35289 23113 35599 23147
rect 35289 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 35599 23113
rect 35289 23051 35599 23085
rect 35289 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 35599 23051
rect 35289 22989 35599 23023
rect 35289 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 35599 22989
rect 35289 14175 35599 22961
rect 35289 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 35599 14175
rect 35289 14113 35599 14147
rect 35289 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 35599 14113
rect 35289 14051 35599 14085
rect 35289 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 35599 14051
rect 35289 13989 35599 14023
rect 35289 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 35599 13989
rect 35289 5175 35599 13961
rect 35289 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 35599 5175
rect 35289 5113 35599 5147
rect 35289 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 35599 5113
rect 35289 5051 35599 5085
rect 35289 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 35599 5051
rect 35289 4989 35599 5023
rect 35289 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 35599 4989
rect 35289 -560 35599 4961
rect 35289 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 35599 -560
rect 35289 -622 35599 -588
rect 35289 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 35599 -622
rect 35289 -684 35599 -650
rect 35289 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 35599 -684
rect 35289 -746 35599 -712
rect 35289 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 35599 -746
rect 35289 -822 35599 -774
rect 48789 298606 49099 299134
rect 48789 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 49099 298606
rect 48789 298544 49099 298578
rect 48789 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 49099 298544
rect 48789 298482 49099 298516
rect 48789 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 49099 298482
rect 48789 298420 49099 298454
rect 48789 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 49099 298420
rect 48789 290175 49099 298392
rect 48789 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 49099 290175
rect 48789 290113 49099 290147
rect 48789 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 49099 290113
rect 48789 290051 49099 290085
rect 48789 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 49099 290051
rect 48789 289989 49099 290023
rect 48789 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 49099 289989
rect 48789 281175 49099 289961
rect 48789 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 49099 281175
rect 48789 281113 49099 281147
rect 48789 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 49099 281113
rect 48789 281051 49099 281085
rect 48789 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 49099 281051
rect 48789 280989 49099 281023
rect 48789 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 49099 280989
rect 48789 272175 49099 280961
rect 48789 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 49099 272175
rect 48789 272113 49099 272147
rect 48789 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 49099 272113
rect 48789 272051 49099 272085
rect 48789 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 49099 272051
rect 48789 271989 49099 272023
rect 48789 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 49099 271989
rect 48789 263175 49099 271961
rect 48789 263147 48837 263175
rect 48865 263147 48899 263175
rect 48927 263147 48961 263175
rect 48989 263147 49023 263175
rect 49051 263147 49099 263175
rect 48789 263113 49099 263147
rect 48789 263085 48837 263113
rect 48865 263085 48899 263113
rect 48927 263085 48961 263113
rect 48989 263085 49023 263113
rect 49051 263085 49099 263113
rect 48789 263051 49099 263085
rect 48789 263023 48837 263051
rect 48865 263023 48899 263051
rect 48927 263023 48961 263051
rect 48989 263023 49023 263051
rect 49051 263023 49099 263051
rect 48789 262989 49099 263023
rect 48789 262961 48837 262989
rect 48865 262961 48899 262989
rect 48927 262961 48961 262989
rect 48989 262961 49023 262989
rect 49051 262961 49099 262989
rect 48789 254175 49099 262961
rect 48789 254147 48837 254175
rect 48865 254147 48899 254175
rect 48927 254147 48961 254175
rect 48989 254147 49023 254175
rect 49051 254147 49099 254175
rect 48789 254113 49099 254147
rect 48789 254085 48837 254113
rect 48865 254085 48899 254113
rect 48927 254085 48961 254113
rect 48989 254085 49023 254113
rect 49051 254085 49099 254113
rect 48789 254051 49099 254085
rect 48789 254023 48837 254051
rect 48865 254023 48899 254051
rect 48927 254023 48961 254051
rect 48989 254023 49023 254051
rect 49051 254023 49099 254051
rect 48789 253989 49099 254023
rect 48789 253961 48837 253989
rect 48865 253961 48899 253989
rect 48927 253961 48961 253989
rect 48989 253961 49023 253989
rect 49051 253961 49099 253989
rect 48789 245175 49099 253961
rect 48789 245147 48837 245175
rect 48865 245147 48899 245175
rect 48927 245147 48961 245175
rect 48989 245147 49023 245175
rect 49051 245147 49099 245175
rect 48789 245113 49099 245147
rect 48789 245085 48837 245113
rect 48865 245085 48899 245113
rect 48927 245085 48961 245113
rect 48989 245085 49023 245113
rect 49051 245085 49099 245113
rect 48789 245051 49099 245085
rect 48789 245023 48837 245051
rect 48865 245023 48899 245051
rect 48927 245023 48961 245051
rect 48989 245023 49023 245051
rect 49051 245023 49099 245051
rect 48789 244989 49099 245023
rect 48789 244961 48837 244989
rect 48865 244961 48899 244989
rect 48927 244961 48961 244989
rect 48989 244961 49023 244989
rect 49051 244961 49099 244989
rect 48789 236175 49099 244961
rect 48789 236147 48837 236175
rect 48865 236147 48899 236175
rect 48927 236147 48961 236175
rect 48989 236147 49023 236175
rect 49051 236147 49099 236175
rect 48789 236113 49099 236147
rect 48789 236085 48837 236113
rect 48865 236085 48899 236113
rect 48927 236085 48961 236113
rect 48989 236085 49023 236113
rect 49051 236085 49099 236113
rect 48789 236051 49099 236085
rect 48789 236023 48837 236051
rect 48865 236023 48899 236051
rect 48927 236023 48961 236051
rect 48989 236023 49023 236051
rect 49051 236023 49099 236051
rect 48789 235989 49099 236023
rect 48789 235961 48837 235989
rect 48865 235961 48899 235989
rect 48927 235961 48961 235989
rect 48989 235961 49023 235989
rect 49051 235961 49099 235989
rect 48789 227175 49099 235961
rect 48789 227147 48837 227175
rect 48865 227147 48899 227175
rect 48927 227147 48961 227175
rect 48989 227147 49023 227175
rect 49051 227147 49099 227175
rect 48789 227113 49099 227147
rect 48789 227085 48837 227113
rect 48865 227085 48899 227113
rect 48927 227085 48961 227113
rect 48989 227085 49023 227113
rect 49051 227085 49099 227113
rect 48789 227051 49099 227085
rect 48789 227023 48837 227051
rect 48865 227023 48899 227051
rect 48927 227023 48961 227051
rect 48989 227023 49023 227051
rect 49051 227023 49099 227051
rect 48789 226989 49099 227023
rect 48789 226961 48837 226989
rect 48865 226961 48899 226989
rect 48927 226961 48961 226989
rect 48989 226961 49023 226989
rect 49051 226961 49099 226989
rect 48789 218175 49099 226961
rect 48789 218147 48837 218175
rect 48865 218147 48899 218175
rect 48927 218147 48961 218175
rect 48989 218147 49023 218175
rect 49051 218147 49099 218175
rect 48789 218113 49099 218147
rect 48789 218085 48837 218113
rect 48865 218085 48899 218113
rect 48927 218085 48961 218113
rect 48989 218085 49023 218113
rect 49051 218085 49099 218113
rect 48789 218051 49099 218085
rect 48789 218023 48837 218051
rect 48865 218023 48899 218051
rect 48927 218023 48961 218051
rect 48989 218023 49023 218051
rect 49051 218023 49099 218051
rect 48789 217989 49099 218023
rect 48789 217961 48837 217989
rect 48865 217961 48899 217989
rect 48927 217961 48961 217989
rect 48989 217961 49023 217989
rect 49051 217961 49099 217989
rect 48789 209175 49099 217961
rect 48789 209147 48837 209175
rect 48865 209147 48899 209175
rect 48927 209147 48961 209175
rect 48989 209147 49023 209175
rect 49051 209147 49099 209175
rect 48789 209113 49099 209147
rect 48789 209085 48837 209113
rect 48865 209085 48899 209113
rect 48927 209085 48961 209113
rect 48989 209085 49023 209113
rect 49051 209085 49099 209113
rect 48789 209051 49099 209085
rect 48789 209023 48837 209051
rect 48865 209023 48899 209051
rect 48927 209023 48961 209051
rect 48989 209023 49023 209051
rect 49051 209023 49099 209051
rect 48789 208989 49099 209023
rect 48789 208961 48837 208989
rect 48865 208961 48899 208989
rect 48927 208961 48961 208989
rect 48989 208961 49023 208989
rect 49051 208961 49099 208989
rect 48789 200175 49099 208961
rect 48789 200147 48837 200175
rect 48865 200147 48899 200175
rect 48927 200147 48961 200175
rect 48989 200147 49023 200175
rect 49051 200147 49099 200175
rect 48789 200113 49099 200147
rect 48789 200085 48837 200113
rect 48865 200085 48899 200113
rect 48927 200085 48961 200113
rect 48989 200085 49023 200113
rect 49051 200085 49099 200113
rect 48789 200051 49099 200085
rect 48789 200023 48837 200051
rect 48865 200023 48899 200051
rect 48927 200023 48961 200051
rect 48989 200023 49023 200051
rect 49051 200023 49099 200051
rect 48789 199989 49099 200023
rect 48789 199961 48837 199989
rect 48865 199961 48899 199989
rect 48927 199961 48961 199989
rect 48989 199961 49023 199989
rect 49051 199961 49099 199989
rect 48789 191175 49099 199961
rect 48789 191147 48837 191175
rect 48865 191147 48899 191175
rect 48927 191147 48961 191175
rect 48989 191147 49023 191175
rect 49051 191147 49099 191175
rect 48789 191113 49099 191147
rect 48789 191085 48837 191113
rect 48865 191085 48899 191113
rect 48927 191085 48961 191113
rect 48989 191085 49023 191113
rect 49051 191085 49099 191113
rect 48789 191051 49099 191085
rect 48789 191023 48837 191051
rect 48865 191023 48899 191051
rect 48927 191023 48961 191051
rect 48989 191023 49023 191051
rect 49051 191023 49099 191051
rect 48789 190989 49099 191023
rect 48789 190961 48837 190989
rect 48865 190961 48899 190989
rect 48927 190961 48961 190989
rect 48989 190961 49023 190989
rect 49051 190961 49099 190989
rect 48789 182175 49099 190961
rect 48789 182147 48837 182175
rect 48865 182147 48899 182175
rect 48927 182147 48961 182175
rect 48989 182147 49023 182175
rect 49051 182147 49099 182175
rect 48789 182113 49099 182147
rect 48789 182085 48837 182113
rect 48865 182085 48899 182113
rect 48927 182085 48961 182113
rect 48989 182085 49023 182113
rect 49051 182085 49099 182113
rect 48789 182051 49099 182085
rect 48789 182023 48837 182051
rect 48865 182023 48899 182051
rect 48927 182023 48961 182051
rect 48989 182023 49023 182051
rect 49051 182023 49099 182051
rect 48789 181989 49099 182023
rect 48789 181961 48837 181989
rect 48865 181961 48899 181989
rect 48927 181961 48961 181989
rect 48989 181961 49023 181989
rect 49051 181961 49099 181989
rect 48789 173175 49099 181961
rect 48789 173147 48837 173175
rect 48865 173147 48899 173175
rect 48927 173147 48961 173175
rect 48989 173147 49023 173175
rect 49051 173147 49099 173175
rect 48789 173113 49099 173147
rect 48789 173085 48837 173113
rect 48865 173085 48899 173113
rect 48927 173085 48961 173113
rect 48989 173085 49023 173113
rect 49051 173085 49099 173113
rect 48789 173051 49099 173085
rect 48789 173023 48837 173051
rect 48865 173023 48899 173051
rect 48927 173023 48961 173051
rect 48989 173023 49023 173051
rect 49051 173023 49099 173051
rect 48789 172989 49099 173023
rect 48789 172961 48837 172989
rect 48865 172961 48899 172989
rect 48927 172961 48961 172989
rect 48989 172961 49023 172989
rect 49051 172961 49099 172989
rect 48789 164175 49099 172961
rect 48789 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 49099 164175
rect 48789 164113 49099 164147
rect 48789 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 49099 164113
rect 48789 164051 49099 164085
rect 48789 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 49099 164051
rect 48789 163989 49099 164023
rect 48789 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 49099 163989
rect 48789 155175 49099 163961
rect 48789 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 49099 155175
rect 48789 155113 49099 155147
rect 48789 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 49099 155113
rect 48789 155051 49099 155085
rect 48789 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 49099 155051
rect 48789 154989 49099 155023
rect 48789 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 49099 154989
rect 48789 146175 49099 154961
rect 48789 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 49099 146175
rect 48789 146113 49099 146147
rect 48789 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 49099 146113
rect 48789 146051 49099 146085
rect 48789 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 49099 146051
rect 48789 145989 49099 146023
rect 48789 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 49099 145989
rect 48789 137175 49099 145961
rect 48789 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 49099 137175
rect 48789 137113 49099 137147
rect 48789 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 49099 137113
rect 48789 137051 49099 137085
rect 48789 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 49099 137051
rect 48789 136989 49099 137023
rect 48789 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 49099 136989
rect 48789 128175 49099 136961
rect 48789 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 49099 128175
rect 48789 128113 49099 128147
rect 48789 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 49099 128113
rect 48789 128051 49099 128085
rect 48789 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 49099 128051
rect 48789 127989 49099 128023
rect 48789 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 49099 127989
rect 48789 119175 49099 127961
rect 48789 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 49099 119175
rect 48789 119113 49099 119147
rect 48789 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 49099 119113
rect 48789 119051 49099 119085
rect 48789 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 49099 119051
rect 48789 118989 49099 119023
rect 48789 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 49099 118989
rect 48789 110175 49099 118961
rect 48789 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 49099 110175
rect 48789 110113 49099 110147
rect 48789 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 49099 110113
rect 48789 110051 49099 110085
rect 48789 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 49099 110051
rect 48789 109989 49099 110023
rect 48789 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 49099 109989
rect 48789 101175 49099 109961
rect 48789 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 49099 101175
rect 48789 101113 49099 101147
rect 48789 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 49099 101113
rect 48789 101051 49099 101085
rect 48789 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 49099 101051
rect 48789 100989 49099 101023
rect 48789 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 49099 100989
rect 48789 92175 49099 100961
rect 48789 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 49099 92175
rect 48789 92113 49099 92147
rect 48789 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 49099 92113
rect 48789 92051 49099 92085
rect 48789 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 49099 92051
rect 48789 91989 49099 92023
rect 48789 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 49099 91989
rect 48789 83175 49099 91961
rect 48789 83147 48837 83175
rect 48865 83147 48899 83175
rect 48927 83147 48961 83175
rect 48989 83147 49023 83175
rect 49051 83147 49099 83175
rect 48789 83113 49099 83147
rect 48789 83085 48837 83113
rect 48865 83085 48899 83113
rect 48927 83085 48961 83113
rect 48989 83085 49023 83113
rect 49051 83085 49099 83113
rect 48789 83051 49099 83085
rect 48789 83023 48837 83051
rect 48865 83023 48899 83051
rect 48927 83023 48961 83051
rect 48989 83023 49023 83051
rect 49051 83023 49099 83051
rect 48789 82989 49099 83023
rect 48789 82961 48837 82989
rect 48865 82961 48899 82989
rect 48927 82961 48961 82989
rect 48989 82961 49023 82989
rect 49051 82961 49099 82989
rect 48789 74175 49099 82961
rect 48789 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 49099 74175
rect 48789 74113 49099 74147
rect 48789 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 49099 74113
rect 48789 74051 49099 74085
rect 48789 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 49099 74051
rect 48789 73989 49099 74023
rect 48789 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 49099 73989
rect 48789 65175 49099 73961
rect 48789 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 49099 65175
rect 48789 65113 49099 65147
rect 48789 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 49099 65113
rect 48789 65051 49099 65085
rect 48789 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 49099 65051
rect 48789 64989 49099 65023
rect 48789 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 49099 64989
rect 48789 56175 49099 64961
rect 48789 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 49099 56175
rect 48789 56113 49099 56147
rect 48789 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 49099 56113
rect 48789 56051 49099 56085
rect 48789 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 49099 56051
rect 48789 55989 49099 56023
rect 48789 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 49099 55989
rect 48789 47175 49099 55961
rect 48789 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 49099 47175
rect 48789 47113 49099 47147
rect 48789 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 49099 47113
rect 48789 47051 49099 47085
rect 48789 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 49099 47051
rect 48789 46989 49099 47023
rect 48789 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 49099 46989
rect 48789 38175 49099 46961
rect 48789 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 49099 38175
rect 48789 38113 49099 38147
rect 48789 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 49099 38113
rect 48789 38051 49099 38085
rect 48789 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 49099 38051
rect 48789 37989 49099 38023
rect 48789 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 49099 37989
rect 48789 29175 49099 37961
rect 48789 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 49099 29175
rect 48789 29113 49099 29147
rect 48789 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 49099 29113
rect 48789 29051 49099 29085
rect 48789 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 49099 29051
rect 48789 28989 49099 29023
rect 48789 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 49099 28989
rect 48789 20175 49099 28961
rect 48789 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 49099 20175
rect 48789 20113 49099 20147
rect 48789 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 49099 20113
rect 48789 20051 49099 20085
rect 48789 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 49099 20051
rect 48789 19989 49099 20023
rect 48789 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 49099 19989
rect 48789 11175 49099 19961
rect 48789 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 49099 11175
rect 48789 11113 49099 11147
rect 48789 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 49099 11113
rect 48789 11051 49099 11085
rect 48789 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 49099 11051
rect 48789 10989 49099 11023
rect 48789 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 49099 10989
rect 48789 2175 49099 10961
rect 48789 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 49099 2175
rect 48789 2113 49099 2147
rect 48789 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 49099 2113
rect 48789 2051 49099 2085
rect 48789 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 49099 2051
rect 48789 1989 49099 2023
rect 48789 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 49099 1989
rect 48789 -80 49099 1961
rect 48789 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 49099 -80
rect 48789 -142 49099 -108
rect 48789 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 49099 -142
rect 48789 -204 49099 -170
rect 48789 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 49099 -204
rect 48789 -266 49099 -232
rect 48789 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 49099 -266
rect 48789 -822 49099 -294
rect 50649 299086 50959 299134
rect 50649 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 50959 299086
rect 50649 299024 50959 299058
rect 50649 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 50959 299024
rect 50649 298962 50959 298996
rect 50649 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 50959 298962
rect 50649 298900 50959 298934
rect 50649 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 50959 298900
rect 50649 293175 50959 298872
rect 50649 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 50959 293175
rect 50649 293113 50959 293147
rect 50649 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 50959 293113
rect 50649 293051 50959 293085
rect 50649 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 50959 293051
rect 50649 292989 50959 293023
rect 50649 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 50959 292989
rect 50649 284175 50959 292961
rect 50649 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 50959 284175
rect 50649 284113 50959 284147
rect 50649 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 50959 284113
rect 50649 284051 50959 284085
rect 50649 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 50959 284051
rect 50649 283989 50959 284023
rect 50649 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 50959 283989
rect 50649 275175 50959 283961
rect 50649 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 50959 275175
rect 50649 275113 50959 275147
rect 50649 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 50959 275113
rect 50649 275051 50959 275085
rect 50649 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 50959 275051
rect 50649 274989 50959 275023
rect 50649 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 50959 274989
rect 50649 266175 50959 274961
rect 50649 266147 50697 266175
rect 50725 266147 50759 266175
rect 50787 266147 50821 266175
rect 50849 266147 50883 266175
rect 50911 266147 50959 266175
rect 50649 266113 50959 266147
rect 50649 266085 50697 266113
rect 50725 266085 50759 266113
rect 50787 266085 50821 266113
rect 50849 266085 50883 266113
rect 50911 266085 50959 266113
rect 50649 266051 50959 266085
rect 50649 266023 50697 266051
rect 50725 266023 50759 266051
rect 50787 266023 50821 266051
rect 50849 266023 50883 266051
rect 50911 266023 50959 266051
rect 50649 265989 50959 266023
rect 50649 265961 50697 265989
rect 50725 265961 50759 265989
rect 50787 265961 50821 265989
rect 50849 265961 50883 265989
rect 50911 265961 50959 265989
rect 50649 257175 50959 265961
rect 50649 257147 50697 257175
rect 50725 257147 50759 257175
rect 50787 257147 50821 257175
rect 50849 257147 50883 257175
rect 50911 257147 50959 257175
rect 50649 257113 50959 257147
rect 50649 257085 50697 257113
rect 50725 257085 50759 257113
rect 50787 257085 50821 257113
rect 50849 257085 50883 257113
rect 50911 257085 50959 257113
rect 50649 257051 50959 257085
rect 50649 257023 50697 257051
rect 50725 257023 50759 257051
rect 50787 257023 50821 257051
rect 50849 257023 50883 257051
rect 50911 257023 50959 257051
rect 50649 256989 50959 257023
rect 50649 256961 50697 256989
rect 50725 256961 50759 256989
rect 50787 256961 50821 256989
rect 50849 256961 50883 256989
rect 50911 256961 50959 256989
rect 50649 248175 50959 256961
rect 50649 248147 50697 248175
rect 50725 248147 50759 248175
rect 50787 248147 50821 248175
rect 50849 248147 50883 248175
rect 50911 248147 50959 248175
rect 50649 248113 50959 248147
rect 50649 248085 50697 248113
rect 50725 248085 50759 248113
rect 50787 248085 50821 248113
rect 50849 248085 50883 248113
rect 50911 248085 50959 248113
rect 50649 248051 50959 248085
rect 50649 248023 50697 248051
rect 50725 248023 50759 248051
rect 50787 248023 50821 248051
rect 50849 248023 50883 248051
rect 50911 248023 50959 248051
rect 50649 247989 50959 248023
rect 50649 247961 50697 247989
rect 50725 247961 50759 247989
rect 50787 247961 50821 247989
rect 50849 247961 50883 247989
rect 50911 247961 50959 247989
rect 50649 239175 50959 247961
rect 50649 239147 50697 239175
rect 50725 239147 50759 239175
rect 50787 239147 50821 239175
rect 50849 239147 50883 239175
rect 50911 239147 50959 239175
rect 50649 239113 50959 239147
rect 50649 239085 50697 239113
rect 50725 239085 50759 239113
rect 50787 239085 50821 239113
rect 50849 239085 50883 239113
rect 50911 239085 50959 239113
rect 50649 239051 50959 239085
rect 50649 239023 50697 239051
rect 50725 239023 50759 239051
rect 50787 239023 50821 239051
rect 50849 239023 50883 239051
rect 50911 239023 50959 239051
rect 50649 238989 50959 239023
rect 50649 238961 50697 238989
rect 50725 238961 50759 238989
rect 50787 238961 50821 238989
rect 50849 238961 50883 238989
rect 50911 238961 50959 238989
rect 50649 230175 50959 238961
rect 50649 230147 50697 230175
rect 50725 230147 50759 230175
rect 50787 230147 50821 230175
rect 50849 230147 50883 230175
rect 50911 230147 50959 230175
rect 50649 230113 50959 230147
rect 50649 230085 50697 230113
rect 50725 230085 50759 230113
rect 50787 230085 50821 230113
rect 50849 230085 50883 230113
rect 50911 230085 50959 230113
rect 50649 230051 50959 230085
rect 50649 230023 50697 230051
rect 50725 230023 50759 230051
rect 50787 230023 50821 230051
rect 50849 230023 50883 230051
rect 50911 230023 50959 230051
rect 50649 229989 50959 230023
rect 50649 229961 50697 229989
rect 50725 229961 50759 229989
rect 50787 229961 50821 229989
rect 50849 229961 50883 229989
rect 50911 229961 50959 229989
rect 50649 221175 50959 229961
rect 50649 221147 50697 221175
rect 50725 221147 50759 221175
rect 50787 221147 50821 221175
rect 50849 221147 50883 221175
rect 50911 221147 50959 221175
rect 50649 221113 50959 221147
rect 50649 221085 50697 221113
rect 50725 221085 50759 221113
rect 50787 221085 50821 221113
rect 50849 221085 50883 221113
rect 50911 221085 50959 221113
rect 50649 221051 50959 221085
rect 50649 221023 50697 221051
rect 50725 221023 50759 221051
rect 50787 221023 50821 221051
rect 50849 221023 50883 221051
rect 50911 221023 50959 221051
rect 50649 220989 50959 221023
rect 50649 220961 50697 220989
rect 50725 220961 50759 220989
rect 50787 220961 50821 220989
rect 50849 220961 50883 220989
rect 50911 220961 50959 220989
rect 50649 212175 50959 220961
rect 50649 212147 50697 212175
rect 50725 212147 50759 212175
rect 50787 212147 50821 212175
rect 50849 212147 50883 212175
rect 50911 212147 50959 212175
rect 50649 212113 50959 212147
rect 50649 212085 50697 212113
rect 50725 212085 50759 212113
rect 50787 212085 50821 212113
rect 50849 212085 50883 212113
rect 50911 212085 50959 212113
rect 50649 212051 50959 212085
rect 50649 212023 50697 212051
rect 50725 212023 50759 212051
rect 50787 212023 50821 212051
rect 50849 212023 50883 212051
rect 50911 212023 50959 212051
rect 50649 211989 50959 212023
rect 50649 211961 50697 211989
rect 50725 211961 50759 211989
rect 50787 211961 50821 211989
rect 50849 211961 50883 211989
rect 50911 211961 50959 211989
rect 50649 203175 50959 211961
rect 50649 203147 50697 203175
rect 50725 203147 50759 203175
rect 50787 203147 50821 203175
rect 50849 203147 50883 203175
rect 50911 203147 50959 203175
rect 50649 203113 50959 203147
rect 50649 203085 50697 203113
rect 50725 203085 50759 203113
rect 50787 203085 50821 203113
rect 50849 203085 50883 203113
rect 50911 203085 50959 203113
rect 50649 203051 50959 203085
rect 50649 203023 50697 203051
rect 50725 203023 50759 203051
rect 50787 203023 50821 203051
rect 50849 203023 50883 203051
rect 50911 203023 50959 203051
rect 50649 202989 50959 203023
rect 50649 202961 50697 202989
rect 50725 202961 50759 202989
rect 50787 202961 50821 202989
rect 50849 202961 50883 202989
rect 50911 202961 50959 202989
rect 50649 194175 50959 202961
rect 50649 194147 50697 194175
rect 50725 194147 50759 194175
rect 50787 194147 50821 194175
rect 50849 194147 50883 194175
rect 50911 194147 50959 194175
rect 50649 194113 50959 194147
rect 50649 194085 50697 194113
rect 50725 194085 50759 194113
rect 50787 194085 50821 194113
rect 50849 194085 50883 194113
rect 50911 194085 50959 194113
rect 50649 194051 50959 194085
rect 50649 194023 50697 194051
rect 50725 194023 50759 194051
rect 50787 194023 50821 194051
rect 50849 194023 50883 194051
rect 50911 194023 50959 194051
rect 50649 193989 50959 194023
rect 50649 193961 50697 193989
rect 50725 193961 50759 193989
rect 50787 193961 50821 193989
rect 50849 193961 50883 193989
rect 50911 193961 50959 193989
rect 50649 185175 50959 193961
rect 50649 185147 50697 185175
rect 50725 185147 50759 185175
rect 50787 185147 50821 185175
rect 50849 185147 50883 185175
rect 50911 185147 50959 185175
rect 50649 185113 50959 185147
rect 50649 185085 50697 185113
rect 50725 185085 50759 185113
rect 50787 185085 50821 185113
rect 50849 185085 50883 185113
rect 50911 185085 50959 185113
rect 50649 185051 50959 185085
rect 50649 185023 50697 185051
rect 50725 185023 50759 185051
rect 50787 185023 50821 185051
rect 50849 185023 50883 185051
rect 50911 185023 50959 185051
rect 50649 184989 50959 185023
rect 50649 184961 50697 184989
rect 50725 184961 50759 184989
rect 50787 184961 50821 184989
rect 50849 184961 50883 184989
rect 50911 184961 50959 184989
rect 50649 176175 50959 184961
rect 50649 176147 50697 176175
rect 50725 176147 50759 176175
rect 50787 176147 50821 176175
rect 50849 176147 50883 176175
rect 50911 176147 50959 176175
rect 50649 176113 50959 176147
rect 50649 176085 50697 176113
rect 50725 176085 50759 176113
rect 50787 176085 50821 176113
rect 50849 176085 50883 176113
rect 50911 176085 50959 176113
rect 50649 176051 50959 176085
rect 50649 176023 50697 176051
rect 50725 176023 50759 176051
rect 50787 176023 50821 176051
rect 50849 176023 50883 176051
rect 50911 176023 50959 176051
rect 50649 175989 50959 176023
rect 50649 175961 50697 175989
rect 50725 175961 50759 175989
rect 50787 175961 50821 175989
rect 50849 175961 50883 175989
rect 50911 175961 50959 175989
rect 50649 167175 50959 175961
rect 50649 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 50959 167175
rect 50649 167113 50959 167147
rect 50649 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 50959 167113
rect 50649 167051 50959 167085
rect 50649 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 50959 167051
rect 50649 166989 50959 167023
rect 50649 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 50959 166989
rect 50649 158175 50959 166961
rect 50649 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 50959 158175
rect 50649 158113 50959 158147
rect 50649 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 50959 158113
rect 50649 158051 50959 158085
rect 50649 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 50959 158051
rect 50649 157989 50959 158023
rect 50649 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 50959 157989
rect 50649 149175 50959 157961
rect 50649 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 50959 149175
rect 50649 149113 50959 149147
rect 50649 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 50959 149113
rect 50649 149051 50959 149085
rect 50649 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 50959 149051
rect 50649 148989 50959 149023
rect 50649 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 50959 148989
rect 50649 140175 50959 148961
rect 50649 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 50959 140175
rect 50649 140113 50959 140147
rect 50649 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 50959 140113
rect 50649 140051 50959 140085
rect 50649 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 50959 140051
rect 50649 139989 50959 140023
rect 50649 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 50959 139989
rect 50649 131175 50959 139961
rect 50649 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 50959 131175
rect 50649 131113 50959 131147
rect 50649 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 50959 131113
rect 50649 131051 50959 131085
rect 50649 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 50959 131051
rect 50649 130989 50959 131023
rect 50649 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 50959 130989
rect 50649 122175 50959 130961
rect 50649 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 50959 122175
rect 50649 122113 50959 122147
rect 50649 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 50959 122113
rect 50649 122051 50959 122085
rect 50649 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 50959 122051
rect 50649 121989 50959 122023
rect 50649 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 50959 121989
rect 50649 113175 50959 121961
rect 50649 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 50959 113175
rect 50649 113113 50959 113147
rect 50649 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 50959 113113
rect 50649 113051 50959 113085
rect 50649 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 50959 113051
rect 50649 112989 50959 113023
rect 50649 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 50959 112989
rect 50649 104175 50959 112961
rect 50649 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 50959 104175
rect 50649 104113 50959 104147
rect 50649 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 50959 104113
rect 50649 104051 50959 104085
rect 50649 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 50959 104051
rect 50649 103989 50959 104023
rect 50649 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 50959 103989
rect 50649 95175 50959 103961
rect 50649 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 50959 95175
rect 50649 95113 50959 95147
rect 50649 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 50959 95113
rect 50649 95051 50959 95085
rect 50649 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 50959 95051
rect 50649 94989 50959 95023
rect 50649 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 50959 94989
rect 50649 86175 50959 94961
rect 50649 86147 50697 86175
rect 50725 86147 50759 86175
rect 50787 86147 50821 86175
rect 50849 86147 50883 86175
rect 50911 86147 50959 86175
rect 50649 86113 50959 86147
rect 50649 86085 50697 86113
rect 50725 86085 50759 86113
rect 50787 86085 50821 86113
rect 50849 86085 50883 86113
rect 50911 86085 50959 86113
rect 50649 86051 50959 86085
rect 50649 86023 50697 86051
rect 50725 86023 50759 86051
rect 50787 86023 50821 86051
rect 50849 86023 50883 86051
rect 50911 86023 50959 86051
rect 50649 85989 50959 86023
rect 50649 85961 50697 85989
rect 50725 85961 50759 85989
rect 50787 85961 50821 85989
rect 50849 85961 50883 85989
rect 50911 85961 50959 85989
rect 50649 77175 50959 85961
rect 50649 77147 50697 77175
rect 50725 77147 50759 77175
rect 50787 77147 50821 77175
rect 50849 77147 50883 77175
rect 50911 77147 50959 77175
rect 50649 77113 50959 77147
rect 50649 77085 50697 77113
rect 50725 77085 50759 77113
rect 50787 77085 50821 77113
rect 50849 77085 50883 77113
rect 50911 77085 50959 77113
rect 50649 77051 50959 77085
rect 50649 77023 50697 77051
rect 50725 77023 50759 77051
rect 50787 77023 50821 77051
rect 50849 77023 50883 77051
rect 50911 77023 50959 77051
rect 50649 76989 50959 77023
rect 50649 76961 50697 76989
rect 50725 76961 50759 76989
rect 50787 76961 50821 76989
rect 50849 76961 50883 76989
rect 50911 76961 50959 76989
rect 50649 68175 50959 76961
rect 50649 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 50959 68175
rect 50649 68113 50959 68147
rect 50649 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 50959 68113
rect 50649 68051 50959 68085
rect 50649 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 50959 68051
rect 50649 67989 50959 68023
rect 50649 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 50959 67989
rect 50649 59175 50959 67961
rect 50649 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 50959 59175
rect 50649 59113 50959 59147
rect 50649 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 50959 59113
rect 50649 59051 50959 59085
rect 50649 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 50959 59051
rect 50649 58989 50959 59023
rect 50649 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 50959 58989
rect 50649 50175 50959 58961
rect 50649 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 50959 50175
rect 50649 50113 50959 50147
rect 50649 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 50959 50113
rect 50649 50051 50959 50085
rect 50649 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 50959 50051
rect 50649 49989 50959 50023
rect 50649 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 50959 49989
rect 50649 41175 50959 49961
rect 50649 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 50959 41175
rect 50649 41113 50959 41147
rect 50649 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 50959 41113
rect 50649 41051 50959 41085
rect 50649 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 50959 41051
rect 50649 40989 50959 41023
rect 50649 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 50959 40989
rect 50649 32175 50959 40961
rect 50649 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 50959 32175
rect 50649 32113 50959 32147
rect 50649 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 50959 32113
rect 50649 32051 50959 32085
rect 50649 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 50959 32051
rect 50649 31989 50959 32023
rect 50649 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 50959 31989
rect 50649 23175 50959 31961
rect 50649 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 50959 23175
rect 50649 23113 50959 23147
rect 50649 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 50959 23113
rect 50649 23051 50959 23085
rect 50649 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 50959 23051
rect 50649 22989 50959 23023
rect 50649 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 50959 22989
rect 50649 14175 50959 22961
rect 50649 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 50959 14175
rect 50649 14113 50959 14147
rect 50649 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 50959 14113
rect 50649 14051 50959 14085
rect 50649 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 50959 14051
rect 50649 13989 50959 14023
rect 50649 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 50959 13989
rect 50649 5175 50959 13961
rect 50649 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 50959 5175
rect 50649 5113 50959 5147
rect 50649 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 50959 5113
rect 50649 5051 50959 5085
rect 50649 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 50959 5051
rect 50649 4989 50959 5023
rect 50649 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 50959 4989
rect 50649 -560 50959 4961
rect 50649 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 50959 -560
rect 50649 -622 50959 -588
rect 50649 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 50959 -622
rect 50649 -684 50959 -650
rect 50649 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 50959 -684
rect 50649 -746 50959 -712
rect 50649 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 50959 -746
rect 50649 -822 50959 -774
rect 64149 298606 64459 299134
rect 64149 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 64459 298606
rect 64149 298544 64459 298578
rect 64149 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 64459 298544
rect 64149 298482 64459 298516
rect 64149 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 64459 298482
rect 64149 298420 64459 298454
rect 64149 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 64459 298420
rect 64149 290175 64459 298392
rect 64149 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 64459 290175
rect 64149 290113 64459 290147
rect 64149 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 64459 290113
rect 64149 290051 64459 290085
rect 64149 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 64459 290051
rect 64149 289989 64459 290023
rect 64149 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 64459 289989
rect 64149 281175 64459 289961
rect 64149 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 64459 281175
rect 64149 281113 64459 281147
rect 64149 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 64459 281113
rect 64149 281051 64459 281085
rect 64149 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 64459 281051
rect 64149 280989 64459 281023
rect 64149 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 64459 280989
rect 64149 272175 64459 280961
rect 64149 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 64459 272175
rect 64149 272113 64459 272147
rect 64149 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 64459 272113
rect 64149 272051 64459 272085
rect 64149 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 64459 272051
rect 64149 271989 64459 272023
rect 64149 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 64459 271989
rect 64149 263175 64459 271961
rect 64149 263147 64197 263175
rect 64225 263147 64259 263175
rect 64287 263147 64321 263175
rect 64349 263147 64383 263175
rect 64411 263147 64459 263175
rect 64149 263113 64459 263147
rect 64149 263085 64197 263113
rect 64225 263085 64259 263113
rect 64287 263085 64321 263113
rect 64349 263085 64383 263113
rect 64411 263085 64459 263113
rect 64149 263051 64459 263085
rect 64149 263023 64197 263051
rect 64225 263023 64259 263051
rect 64287 263023 64321 263051
rect 64349 263023 64383 263051
rect 64411 263023 64459 263051
rect 64149 262989 64459 263023
rect 64149 262961 64197 262989
rect 64225 262961 64259 262989
rect 64287 262961 64321 262989
rect 64349 262961 64383 262989
rect 64411 262961 64459 262989
rect 64149 254175 64459 262961
rect 64149 254147 64197 254175
rect 64225 254147 64259 254175
rect 64287 254147 64321 254175
rect 64349 254147 64383 254175
rect 64411 254147 64459 254175
rect 64149 254113 64459 254147
rect 64149 254085 64197 254113
rect 64225 254085 64259 254113
rect 64287 254085 64321 254113
rect 64349 254085 64383 254113
rect 64411 254085 64459 254113
rect 64149 254051 64459 254085
rect 64149 254023 64197 254051
rect 64225 254023 64259 254051
rect 64287 254023 64321 254051
rect 64349 254023 64383 254051
rect 64411 254023 64459 254051
rect 64149 253989 64459 254023
rect 64149 253961 64197 253989
rect 64225 253961 64259 253989
rect 64287 253961 64321 253989
rect 64349 253961 64383 253989
rect 64411 253961 64459 253989
rect 64149 245175 64459 253961
rect 64149 245147 64197 245175
rect 64225 245147 64259 245175
rect 64287 245147 64321 245175
rect 64349 245147 64383 245175
rect 64411 245147 64459 245175
rect 64149 245113 64459 245147
rect 64149 245085 64197 245113
rect 64225 245085 64259 245113
rect 64287 245085 64321 245113
rect 64349 245085 64383 245113
rect 64411 245085 64459 245113
rect 64149 245051 64459 245085
rect 64149 245023 64197 245051
rect 64225 245023 64259 245051
rect 64287 245023 64321 245051
rect 64349 245023 64383 245051
rect 64411 245023 64459 245051
rect 64149 244989 64459 245023
rect 64149 244961 64197 244989
rect 64225 244961 64259 244989
rect 64287 244961 64321 244989
rect 64349 244961 64383 244989
rect 64411 244961 64459 244989
rect 64149 236175 64459 244961
rect 64149 236147 64197 236175
rect 64225 236147 64259 236175
rect 64287 236147 64321 236175
rect 64349 236147 64383 236175
rect 64411 236147 64459 236175
rect 64149 236113 64459 236147
rect 64149 236085 64197 236113
rect 64225 236085 64259 236113
rect 64287 236085 64321 236113
rect 64349 236085 64383 236113
rect 64411 236085 64459 236113
rect 64149 236051 64459 236085
rect 64149 236023 64197 236051
rect 64225 236023 64259 236051
rect 64287 236023 64321 236051
rect 64349 236023 64383 236051
rect 64411 236023 64459 236051
rect 64149 235989 64459 236023
rect 64149 235961 64197 235989
rect 64225 235961 64259 235989
rect 64287 235961 64321 235989
rect 64349 235961 64383 235989
rect 64411 235961 64459 235989
rect 64149 227175 64459 235961
rect 64149 227147 64197 227175
rect 64225 227147 64259 227175
rect 64287 227147 64321 227175
rect 64349 227147 64383 227175
rect 64411 227147 64459 227175
rect 64149 227113 64459 227147
rect 64149 227085 64197 227113
rect 64225 227085 64259 227113
rect 64287 227085 64321 227113
rect 64349 227085 64383 227113
rect 64411 227085 64459 227113
rect 64149 227051 64459 227085
rect 64149 227023 64197 227051
rect 64225 227023 64259 227051
rect 64287 227023 64321 227051
rect 64349 227023 64383 227051
rect 64411 227023 64459 227051
rect 64149 226989 64459 227023
rect 64149 226961 64197 226989
rect 64225 226961 64259 226989
rect 64287 226961 64321 226989
rect 64349 226961 64383 226989
rect 64411 226961 64459 226989
rect 64149 218175 64459 226961
rect 64149 218147 64197 218175
rect 64225 218147 64259 218175
rect 64287 218147 64321 218175
rect 64349 218147 64383 218175
rect 64411 218147 64459 218175
rect 64149 218113 64459 218147
rect 64149 218085 64197 218113
rect 64225 218085 64259 218113
rect 64287 218085 64321 218113
rect 64349 218085 64383 218113
rect 64411 218085 64459 218113
rect 64149 218051 64459 218085
rect 64149 218023 64197 218051
rect 64225 218023 64259 218051
rect 64287 218023 64321 218051
rect 64349 218023 64383 218051
rect 64411 218023 64459 218051
rect 64149 217989 64459 218023
rect 64149 217961 64197 217989
rect 64225 217961 64259 217989
rect 64287 217961 64321 217989
rect 64349 217961 64383 217989
rect 64411 217961 64459 217989
rect 64149 209175 64459 217961
rect 64149 209147 64197 209175
rect 64225 209147 64259 209175
rect 64287 209147 64321 209175
rect 64349 209147 64383 209175
rect 64411 209147 64459 209175
rect 64149 209113 64459 209147
rect 64149 209085 64197 209113
rect 64225 209085 64259 209113
rect 64287 209085 64321 209113
rect 64349 209085 64383 209113
rect 64411 209085 64459 209113
rect 64149 209051 64459 209085
rect 64149 209023 64197 209051
rect 64225 209023 64259 209051
rect 64287 209023 64321 209051
rect 64349 209023 64383 209051
rect 64411 209023 64459 209051
rect 64149 208989 64459 209023
rect 64149 208961 64197 208989
rect 64225 208961 64259 208989
rect 64287 208961 64321 208989
rect 64349 208961 64383 208989
rect 64411 208961 64459 208989
rect 64149 200175 64459 208961
rect 64149 200147 64197 200175
rect 64225 200147 64259 200175
rect 64287 200147 64321 200175
rect 64349 200147 64383 200175
rect 64411 200147 64459 200175
rect 64149 200113 64459 200147
rect 64149 200085 64197 200113
rect 64225 200085 64259 200113
rect 64287 200085 64321 200113
rect 64349 200085 64383 200113
rect 64411 200085 64459 200113
rect 64149 200051 64459 200085
rect 64149 200023 64197 200051
rect 64225 200023 64259 200051
rect 64287 200023 64321 200051
rect 64349 200023 64383 200051
rect 64411 200023 64459 200051
rect 64149 199989 64459 200023
rect 64149 199961 64197 199989
rect 64225 199961 64259 199989
rect 64287 199961 64321 199989
rect 64349 199961 64383 199989
rect 64411 199961 64459 199989
rect 64149 191175 64459 199961
rect 64149 191147 64197 191175
rect 64225 191147 64259 191175
rect 64287 191147 64321 191175
rect 64349 191147 64383 191175
rect 64411 191147 64459 191175
rect 64149 191113 64459 191147
rect 64149 191085 64197 191113
rect 64225 191085 64259 191113
rect 64287 191085 64321 191113
rect 64349 191085 64383 191113
rect 64411 191085 64459 191113
rect 64149 191051 64459 191085
rect 64149 191023 64197 191051
rect 64225 191023 64259 191051
rect 64287 191023 64321 191051
rect 64349 191023 64383 191051
rect 64411 191023 64459 191051
rect 64149 190989 64459 191023
rect 64149 190961 64197 190989
rect 64225 190961 64259 190989
rect 64287 190961 64321 190989
rect 64349 190961 64383 190989
rect 64411 190961 64459 190989
rect 64149 182175 64459 190961
rect 64149 182147 64197 182175
rect 64225 182147 64259 182175
rect 64287 182147 64321 182175
rect 64349 182147 64383 182175
rect 64411 182147 64459 182175
rect 64149 182113 64459 182147
rect 64149 182085 64197 182113
rect 64225 182085 64259 182113
rect 64287 182085 64321 182113
rect 64349 182085 64383 182113
rect 64411 182085 64459 182113
rect 64149 182051 64459 182085
rect 64149 182023 64197 182051
rect 64225 182023 64259 182051
rect 64287 182023 64321 182051
rect 64349 182023 64383 182051
rect 64411 182023 64459 182051
rect 64149 181989 64459 182023
rect 64149 181961 64197 181989
rect 64225 181961 64259 181989
rect 64287 181961 64321 181989
rect 64349 181961 64383 181989
rect 64411 181961 64459 181989
rect 64149 173175 64459 181961
rect 64149 173147 64197 173175
rect 64225 173147 64259 173175
rect 64287 173147 64321 173175
rect 64349 173147 64383 173175
rect 64411 173147 64459 173175
rect 64149 173113 64459 173147
rect 64149 173085 64197 173113
rect 64225 173085 64259 173113
rect 64287 173085 64321 173113
rect 64349 173085 64383 173113
rect 64411 173085 64459 173113
rect 64149 173051 64459 173085
rect 64149 173023 64197 173051
rect 64225 173023 64259 173051
rect 64287 173023 64321 173051
rect 64349 173023 64383 173051
rect 64411 173023 64459 173051
rect 64149 172989 64459 173023
rect 64149 172961 64197 172989
rect 64225 172961 64259 172989
rect 64287 172961 64321 172989
rect 64349 172961 64383 172989
rect 64411 172961 64459 172989
rect 64149 164175 64459 172961
rect 64149 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 64459 164175
rect 64149 164113 64459 164147
rect 64149 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 64459 164113
rect 64149 164051 64459 164085
rect 64149 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 64459 164051
rect 64149 163989 64459 164023
rect 64149 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 64459 163989
rect 64149 155175 64459 163961
rect 64149 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 64459 155175
rect 64149 155113 64459 155147
rect 64149 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 64459 155113
rect 64149 155051 64459 155085
rect 64149 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 64459 155051
rect 64149 154989 64459 155023
rect 64149 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 64459 154989
rect 64149 146175 64459 154961
rect 64149 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 64459 146175
rect 64149 146113 64459 146147
rect 64149 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 64459 146113
rect 64149 146051 64459 146085
rect 64149 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 64459 146051
rect 64149 145989 64459 146023
rect 64149 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 64459 145989
rect 64149 137175 64459 145961
rect 64149 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 64459 137175
rect 64149 137113 64459 137147
rect 64149 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 64459 137113
rect 64149 137051 64459 137085
rect 64149 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 64459 137051
rect 64149 136989 64459 137023
rect 64149 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 64459 136989
rect 64149 128175 64459 136961
rect 64149 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 64459 128175
rect 64149 128113 64459 128147
rect 64149 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 64459 128113
rect 64149 128051 64459 128085
rect 64149 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 64459 128051
rect 64149 127989 64459 128023
rect 64149 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 64459 127989
rect 64149 119175 64459 127961
rect 64149 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 64459 119175
rect 64149 119113 64459 119147
rect 64149 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 64459 119113
rect 64149 119051 64459 119085
rect 64149 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 64459 119051
rect 64149 118989 64459 119023
rect 64149 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 64459 118989
rect 64149 110175 64459 118961
rect 64149 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 64459 110175
rect 64149 110113 64459 110147
rect 64149 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 64459 110113
rect 64149 110051 64459 110085
rect 64149 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 64459 110051
rect 64149 109989 64459 110023
rect 64149 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 64459 109989
rect 64149 101175 64459 109961
rect 64149 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 64459 101175
rect 64149 101113 64459 101147
rect 64149 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 64459 101113
rect 64149 101051 64459 101085
rect 64149 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 64459 101051
rect 64149 100989 64459 101023
rect 64149 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 64459 100989
rect 64149 92175 64459 100961
rect 64149 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 64459 92175
rect 64149 92113 64459 92147
rect 64149 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 64459 92113
rect 64149 92051 64459 92085
rect 64149 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 64459 92051
rect 64149 91989 64459 92023
rect 64149 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 64459 91989
rect 64149 83175 64459 91961
rect 64149 83147 64197 83175
rect 64225 83147 64259 83175
rect 64287 83147 64321 83175
rect 64349 83147 64383 83175
rect 64411 83147 64459 83175
rect 64149 83113 64459 83147
rect 64149 83085 64197 83113
rect 64225 83085 64259 83113
rect 64287 83085 64321 83113
rect 64349 83085 64383 83113
rect 64411 83085 64459 83113
rect 64149 83051 64459 83085
rect 64149 83023 64197 83051
rect 64225 83023 64259 83051
rect 64287 83023 64321 83051
rect 64349 83023 64383 83051
rect 64411 83023 64459 83051
rect 64149 82989 64459 83023
rect 64149 82961 64197 82989
rect 64225 82961 64259 82989
rect 64287 82961 64321 82989
rect 64349 82961 64383 82989
rect 64411 82961 64459 82989
rect 64149 74175 64459 82961
rect 64149 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 64459 74175
rect 64149 74113 64459 74147
rect 64149 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 64459 74113
rect 64149 74051 64459 74085
rect 64149 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 64459 74051
rect 64149 73989 64459 74023
rect 64149 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 64459 73989
rect 64149 65175 64459 73961
rect 64149 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 64459 65175
rect 64149 65113 64459 65147
rect 64149 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 64459 65113
rect 64149 65051 64459 65085
rect 64149 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 64459 65051
rect 64149 64989 64459 65023
rect 64149 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 64459 64989
rect 64149 56175 64459 64961
rect 64149 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 64459 56175
rect 64149 56113 64459 56147
rect 64149 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 64459 56113
rect 64149 56051 64459 56085
rect 64149 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 64459 56051
rect 64149 55989 64459 56023
rect 64149 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 64459 55989
rect 64149 47175 64459 55961
rect 64149 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 64459 47175
rect 64149 47113 64459 47147
rect 64149 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 64459 47113
rect 64149 47051 64459 47085
rect 64149 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 64459 47051
rect 64149 46989 64459 47023
rect 64149 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 64459 46989
rect 64149 38175 64459 46961
rect 64149 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 64459 38175
rect 64149 38113 64459 38147
rect 64149 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 64459 38113
rect 64149 38051 64459 38085
rect 64149 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 64459 38051
rect 64149 37989 64459 38023
rect 64149 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 64459 37989
rect 64149 29175 64459 37961
rect 64149 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 64459 29175
rect 64149 29113 64459 29147
rect 64149 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 64459 29113
rect 64149 29051 64459 29085
rect 64149 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 64459 29051
rect 64149 28989 64459 29023
rect 64149 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 64459 28989
rect 64149 20175 64459 28961
rect 64149 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 64459 20175
rect 64149 20113 64459 20147
rect 64149 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 64459 20113
rect 64149 20051 64459 20085
rect 64149 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 64459 20051
rect 64149 19989 64459 20023
rect 64149 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 64459 19989
rect 64149 11175 64459 19961
rect 64149 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 64459 11175
rect 64149 11113 64459 11147
rect 64149 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 64459 11113
rect 64149 11051 64459 11085
rect 64149 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 64459 11051
rect 64149 10989 64459 11023
rect 64149 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 64459 10989
rect 64149 2175 64459 10961
rect 64149 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 64459 2175
rect 64149 2113 64459 2147
rect 64149 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 64459 2113
rect 64149 2051 64459 2085
rect 64149 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 64459 2051
rect 64149 1989 64459 2023
rect 64149 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 64459 1989
rect 64149 -80 64459 1961
rect 64149 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 64459 -80
rect 64149 -142 64459 -108
rect 64149 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 64459 -142
rect 64149 -204 64459 -170
rect 64149 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 64459 -204
rect 64149 -266 64459 -232
rect 64149 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 64459 -266
rect 64149 -822 64459 -294
rect 66009 299086 66319 299134
rect 66009 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 66319 299086
rect 66009 299024 66319 299058
rect 66009 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 66319 299024
rect 66009 298962 66319 298996
rect 66009 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 66319 298962
rect 66009 298900 66319 298934
rect 66009 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 66319 298900
rect 66009 293175 66319 298872
rect 66009 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 66319 293175
rect 66009 293113 66319 293147
rect 66009 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 66319 293113
rect 66009 293051 66319 293085
rect 66009 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 66319 293051
rect 66009 292989 66319 293023
rect 66009 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 66319 292989
rect 66009 284175 66319 292961
rect 66009 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 66319 284175
rect 66009 284113 66319 284147
rect 66009 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 66319 284113
rect 66009 284051 66319 284085
rect 66009 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 66319 284051
rect 66009 283989 66319 284023
rect 66009 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 66319 283989
rect 66009 275175 66319 283961
rect 66009 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 66319 275175
rect 66009 275113 66319 275147
rect 66009 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 66319 275113
rect 66009 275051 66319 275085
rect 66009 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 66319 275051
rect 66009 274989 66319 275023
rect 66009 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 66319 274989
rect 66009 266175 66319 274961
rect 66009 266147 66057 266175
rect 66085 266147 66119 266175
rect 66147 266147 66181 266175
rect 66209 266147 66243 266175
rect 66271 266147 66319 266175
rect 66009 266113 66319 266147
rect 66009 266085 66057 266113
rect 66085 266085 66119 266113
rect 66147 266085 66181 266113
rect 66209 266085 66243 266113
rect 66271 266085 66319 266113
rect 66009 266051 66319 266085
rect 66009 266023 66057 266051
rect 66085 266023 66119 266051
rect 66147 266023 66181 266051
rect 66209 266023 66243 266051
rect 66271 266023 66319 266051
rect 66009 265989 66319 266023
rect 66009 265961 66057 265989
rect 66085 265961 66119 265989
rect 66147 265961 66181 265989
rect 66209 265961 66243 265989
rect 66271 265961 66319 265989
rect 66009 257175 66319 265961
rect 66009 257147 66057 257175
rect 66085 257147 66119 257175
rect 66147 257147 66181 257175
rect 66209 257147 66243 257175
rect 66271 257147 66319 257175
rect 66009 257113 66319 257147
rect 66009 257085 66057 257113
rect 66085 257085 66119 257113
rect 66147 257085 66181 257113
rect 66209 257085 66243 257113
rect 66271 257085 66319 257113
rect 66009 257051 66319 257085
rect 66009 257023 66057 257051
rect 66085 257023 66119 257051
rect 66147 257023 66181 257051
rect 66209 257023 66243 257051
rect 66271 257023 66319 257051
rect 66009 256989 66319 257023
rect 66009 256961 66057 256989
rect 66085 256961 66119 256989
rect 66147 256961 66181 256989
rect 66209 256961 66243 256989
rect 66271 256961 66319 256989
rect 66009 248175 66319 256961
rect 66009 248147 66057 248175
rect 66085 248147 66119 248175
rect 66147 248147 66181 248175
rect 66209 248147 66243 248175
rect 66271 248147 66319 248175
rect 66009 248113 66319 248147
rect 66009 248085 66057 248113
rect 66085 248085 66119 248113
rect 66147 248085 66181 248113
rect 66209 248085 66243 248113
rect 66271 248085 66319 248113
rect 66009 248051 66319 248085
rect 66009 248023 66057 248051
rect 66085 248023 66119 248051
rect 66147 248023 66181 248051
rect 66209 248023 66243 248051
rect 66271 248023 66319 248051
rect 66009 247989 66319 248023
rect 66009 247961 66057 247989
rect 66085 247961 66119 247989
rect 66147 247961 66181 247989
rect 66209 247961 66243 247989
rect 66271 247961 66319 247989
rect 66009 239175 66319 247961
rect 66009 239147 66057 239175
rect 66085 239147 66119 239175
rect 66147 239147 66181 239175
rect 66209 239147 66243 239175
rect 66271 239147 66319 239175
rect 66009 239113 66319 239147
rect 66009 239085 66057 239113
rect 66085 239085 66119 239113
rect 66147 239085 66181 239113
rect 66209 239085 66243 239113
rect 66271 239085 66319 239113
rect 66009 239051 66319 239085
rect 66009 239023 66057 239051
rect 66085 239023 66119 239051
rect 66147 239023 66181 239051
rect 66209 239023 66243 239051
rect 66271 239023 66319 239051
rect 66009 238989 66319 239023
rect 66009 238961 66057 238989
rect 66085 238961 66119 238989
rect 66147 238961 66181 238989
rect 66209 238961 66243 238989
rect 66271 238961 66319 238989
rect 66009 230175 66319 238961
rect 66009 230147 66057 230175
rect 66085 230147 66119 230175
rect 66147 230147 66181 230175
rect 66209 230147 66243 230175
rect 66271 230147 66319 230175
rect 66009 230113 66319 230147
rect 66009 230085 66057 230113
rect 66085 230085 66119 230113
rect 66147 230085 66181 230113
rect 66209 230085 66243 230113
rect 66271 230085 66319 230113
rect 66009 230051 66319 230085
rect 66009 230023 66057 230051
rect 66085 230023 66119 230051
rect 66147 230023 66181 230051
rect 66209 230023 66243 230051
rect 66271 230023 66319 230051
rect 66009 229989 66319 230023
rect 66009 229961 66057 229989
rect 66085 229961 66119 229989
rect 66147 229961 66181 229989
rect 66209 229961 66243 229989
rect 66271 229961 66319 229989
rect 66009 221175 66319 229961
rect 66009 221147 66057 221175
rect 66085 221147 66119 221175
rect 66147 221147 66181 221175
rect 66209 221147 66243 221175
rect 66271 221147 66319 221175
rect 66009 221113 66319 221147
rect 66009 221085 66057 221113
rect 66085 221085 66119 221113
rect 66147 221085 66181 221113
rect 66209 221085 66243 221113
rect 66271 221085 66319 221113
rect 66009 221051 66319 221085
rect 66009 221023 66057 221051
rect 66085 221023 66119 221051
rect 66147 221023 66181 221051
rect 66209 221023 66243 221051
rect 66271 221023 66319 221051
rect 66009 220989 66319 221023
rect 66009 220961 66057 220989
rect 66085 220961 66119 220989
rect 66147 220961 66181 220989
rect 66209 220961 66243 220989
rect 66271 220961 66319 220989
rect 66009 212175 66319 220961
rect 66009 212147 66057 212175
rect 66085 212147 66119 212175
rect 66147 212147 66181 212175
rect 66209 212147 66243 212175
rect 66271 212147 66319 212175
rect 66009 212113 66319 212147
rect 66009 212085 66057 212113
rect 66085 212085 66119 212113
rect 66147 212085 66181 212113
rect 66209 212085 66243 212113
rect 66271 212085 66319 212113
rect 66009 212051 66319 212085
rect 66009 212023 66057 212051
rect 66085 212023 66119 212051
rect 66147 212023 66181 212051
rect 66209 212023 66243 212051
rect 66271 212023 66319 212051
rect 66009 211989 66319 212023
rect 66009 211961 66057 211989
rect 66085 211961 66119 211989
rect 66147 211961 66181 211989
rect 66209 211961 66243 211989
rect 66271 211961 66319 211989
rect 66009 203175 66319 211961
rect 66009 203147 66057 203175
rect 66085 203147 66119 203175
rect 66147 203147 66181 203175
rect 66209 203147 66243 203175
rect 66271 203147 66319 203175
rect 66009 203113 66319 203147
rect 66009 203085 66057 203113
rect 66085 203085 66119 203113
rect 66147 203085 66181 203113
rect 66209 203085 66243 203113
rect 66271 203085 66319 203113
rect 66009 203051 66319 203085
rect 66009 203023 66057 203051
rect 66085 203023 66119 203051
rect 66147 203023 66181 203051
rect 66209 203023 66243 203051
rect 66271 203023 66319 203051
rect 66009 202989 66319 203023
rect 66009 202961 66057 202989
rect 66085 202961 66119 202989
rect 66147 202961 66181 202989
rect 66209 202961 66243 202989
rect 66271 202961 66319 202989
rect 66009 194175 66319 202961
rect 66009 194147 66057 194175
rect 66085 194147 66119 194175
rect 66147 194147 66181 194175
rect 66209 194147 66243 194175
rect 66271 194147 66319 194175
rect 66009 194113 66319 194147
rect 66009 194085 66057 194113
rect 66085 194085 66119 194113
rect 66147 194085 66181 194113
rect 66209 194085 66243 194113
rect 66271 194085 66319 194113
rect 66009 194051 66319 194085
rect 66009 194023 66057 194051
rect 66085 194023 66119 194051
rect 66147 194023 66181 194051
rect 66209 194023 66243 194051
rect 66271 194023 66319 194051
rect 66009 193989 66319 194023
rect 66009 193961 66057 193989
rect 66085 193961 66119 193989
rect 66147 193961 66181 193989
rect 66209 193961 66243 193989
rect 66271 193961 66319 193989
rect 66009 185175 66319 193961
rect 66009 185147 66057 185175
rect 66085 185147 66119 185175
rect 66147 185147 66181 185175
rect 66209 185147 66243 185175
rect 66271 185147 66319 185175
rect 66009 185113 66319 185147
rect 66009 185085 66057 185113
rect 66085 185085 66119 185113
rect 66147 185085 66181 185113
rect 66209 185085 66243 185113
rect 66271 185085 66319 185113
rect 66009 185051 66319 185085
rect 66009 185023 66057 185051
rect 66085 185023 66119 185051
rect 66147 185023 66181 185051
rect 66209 185023 66243 185051
rect 66271 185023 66319 185051
rect 66009 184989 66319 185023
rect 66009 184961 66057 184989
rect 66085 184961 66119 184989
rect 66147 184961 66181 184989
rect 66209 184961 66243 184989
rect 66271 184961 66319 184989
rect 66009 176175 66319 184961
rect 66009 176147 66057 176175
rect 66085 176147 66119 176175
rect 66147 176147 66181 176175
rect 66209 176147 66243 176175
rect 66271 176147 66319 176175
rect 66009 176113 66319 176147
rect 66009 176085 66057 176113
rect 66085 176085 66119 176113
rect 66147 176085 66181 176113
rect 66209 176085 66243 176113
rect 66271 176085 66319 176113
rect 66009 176051 66319 176085
rect 66009 176023 66057 176051
rect 66085 176023 66119 176051
rect 66147 176023 66181 176051
rect 66209 176023 66243 176051
rect 66271 176023 66319 176051
rect 66009 175989 66319 176023
rect 66009 175961 66057 175989
rect 66085 175961 66119 175989
rect 66147 175961 66181 175989
rect 66209 175961 66243 175989
rect 66271 175961 66319 175989
rect 66009 167175 66319 175961
rect 66009 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 66319 167175
rect 66009 167113 66319 167147
rect 66009 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 66319 167113
rect 66009 167051 66319 167085
rect 66009 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 66319 167051
rect 66009 166989 66319 167023
rect 66009 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 66319 166989
rect 66009 158175 66319 166961
rect 66009 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 66319 158175
rect 66009 158113 66319 158147
rect 66009 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 66319 158113
rect 66009 158051 66319 158085
rect 66009 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 66319 158051
rect 66009 157989 66319 158023
rect 66009 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 66319 157989
rect 66009 149175 66319 157961
rect 66009 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 66319 149175
rect 66009 149113 66319 149147
rect 66009 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 66319 149113
rect 66009 149051 66319 149085
rect 66009 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 66319 149051
rect 66009 148989 66319 149023
rect 66009 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 66319 148989
rect 66009 140175 66319 148961
rect 66009 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 66319 140175
rect 66009 140113 66319 140147
rect 66009 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 66319 140113
rect 66009 140051 66319 140085
rect 66009 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 66319 140051
rect 66009 139989 66319 140023
rect 66009 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 66319 139989
rect 66009 131175 66319 139961
rect 66009 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 66319 131175
rect 66009 131113 66319 131147
rect 66009 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 66319 131113
rect 66009 131051 66319 131085
rect 66009 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 66319 131051
rect 66009 130989 66319 131023
rect 66009 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 66319 130989
rect 66009 122175 66319 130961
rect 66009 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 66319 122175
rect 66009 122113 66319 122147
rect 66009 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 66319 122113
rect 66009 122051 66319 122085
rect 66009 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 66319 122051
rect 66009 121989 66319 122023
rect 66009 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 66319 121989
rect 66009 113175 66319 121961
rect 66009 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 66319 113175
rect 66009 113113 66319 113147
rect 66009 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 66319 113113
rect 66009 113051 66319 113085
rect 66009 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 66319 113051
rect 66009 112989 66319 113023
rect 66009 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 66319 112989
rect 66009 104175 66319 112961
rect 66009 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 66319 104175
rect 66009 104113 66319 104147
rect 66009 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 66319 104113
rect 66009 104051 66319 104085
rect 66009 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 66319 104051
rect 66009 103989 66319 104023
rect 66009 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 66319 103989
rect 66009 95175 66319 103961
rect 66009 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 66319 95175
rect 66009 95113 66319 95147
rect 66009 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 66319 95113
rect 66009 95051 66319 95085
rect 66009 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 66319 95051
rect 66009 94989 66319 95023
rect 66009 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 66319 94989
rect 66009 86175 66319 94961
rect 66009 86147 66057 86175
rect 66085 86147 66119 86175
rect 66147 86147 66181 86175
rect 66209 86147 66243 86175
rect 66271 86147 66319 86175
rect 66009 86113 66319 86147
rect 66009 86085 66057 86113
rect 66085 86085 66119 86113
rect 66147 86085 66181 86113
rect 66209 86085 66243 86113
rect 66271 86085 66319 86113
rect 66009 86051 66319 86085
rect 66009 86023 66057 86051
rect 66085 86023 66119 86051
rect 66147 86023 66181 86051
rect 66209 86023 66243 86051
rect 66271 86023 66319 86051
rect 66009 85989 66319 86023
rect 66009 85961 66057 85989
rect 66085 85961 66119 85989
rect 66147 85961 66181 85989
rect 66209 85961 66243 85989
rect 66271 85961 66319 85989
rect 66009 77175 66319 85961
rect 66009 77147 66057 77175
rect 66085 77147 66119 77175
rect 66147 77147 66181 77175
rect 66209 77147 66243 77175
rect 66271 77147 66319 77175
rect 66009 77113 66319 77147
rect 66009 77085 66057 77113
rect 66085 77085 66119 77113
rect 66147 77085 66181 77113
rect 66209 77085 66243 77113
rect 66271 77085 66319 77113
rect 66009 77051 66319 77085
rect 66009 77023 66057 77051
rect 66085 77023 66119 77051
rect 66147 77023 66181 77051
rect 66209 77023 66243 77051
rect 66271 77023 66319 77051
rect 66009 76989 66319 77023
rect 66009 76961 66057 76989
rect 66085 76961 66119 76989
rect 66147 76961 66181 76989
rect 66209 76961 66243 76989
rect 66271 76961 66319 76989
rect 66009 68175 66319 76961
rect 66009 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 66319 68175
rect 66009 68113 66319 68147
rect 66009 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 66319 68113
rect 66009 68051 66319 68085
rect 66009 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 66319 68051
rect 66009 67989 66319 68023
rect 66009 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 66319 67989
rect 66009 59175 66319 67961
rect 66009 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 66319 59175
rect 66009 59113 66319 59147
rect 66009 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 66319 59113
rect 66009 59051 66319 59085
rect 66009 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 66319 59051
rect 66009 58989 66319 59023
rect 66009 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 66319 58989
rect 66009 50175 66319 58961
rect 66009 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 66319 50175
rect 66009 50113 66319 50147
rect 66009 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 66319 50113
rect 66009 50051 66319 50085
rect 66009 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 66319 50051
rect 66009 49989 66319 50023
rect 66009 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 66319 49989
rect 66009 41175 66319 49961
rect 66009 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 66319 41175
rect 66009 41113 66319 41147
rect 66009 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 66319 41113
rect 66009 41051 66319 41085
rect 66009 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 66319 41051
rect 66009 40989 66319 41023
rect 66009 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 66319 40989
rect 66009 32175 66319 40961
rect 66009 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 66319 32175
rect 66009 32113 66319 32147
rect 66009 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 66319 32113
rect 66009 32051 66319 32085
rect 66009 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 66319 32051
rect 66009 31989 66319 32023
rect 66009 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 66319 31989
rect 66009 23175 66319 31961
rect 66009 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 66319 23175
rect 66009 23113 66319 23147
rect 66009 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 66319 23113
rect 66009 23051 66319 23085
rect 66009 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 66319 23051
rect 66009 22989 66319 23023
rect 66009 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 66319 22989
rect 66009 14175 66319 22961
rect 66009 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 66319 14175
rect 66009 14113 66319 14147
rect 66009 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 66319 14113
rect 66009 14051 66319 14085
rect 66009 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 66319 14051
rect 66009 13989 66319 14023
rect 66009 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 66319 13989
rect 66009 5175 66319 13961
rect 66009 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 66319 5175
rect 66009 5113 66319 5147
rect 66009 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 66319 5113
rect 66009 5051 66319 5085
rect 66009 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 66319 5051
rect 66009 4989 66319 5023
rect 66009 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 66319 4989
rect 66009 -560 66319 4961
rect 66009 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 66319 -560
rect 66009 -622 66319 -588
rect 66009 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 66319 -622
rect 66009 -684 66319 -650
rect 66009 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 66319 -684
rect 66009 -746 66319 -712
rect 66009 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 66319 -746
rect 66009 -822 66319 -774
rect 79509 298606 79819 299134
rect 79509 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 79819 298606
rect 79509 298544 79819 298578
rect 79509 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 79819 298544
rect 79509 298482 79819 298516
rect 79509 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 79819 298482
rect 79509 298420 79819 298454
rect 79509 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 79819 298420
rect 79509 290175 79819 298392
rect 79509 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 79819 290175
rect 79509 290113 79819 290147
rect 79509 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 79819 290113
rect 79509 290051 79819 290085
rect 79509 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 79819 290051
rect 79509 289989 79819 290023
rect 79509 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 79819 289989
rect 79509 281175 79819 289961
rect 79509 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 79819 281175
rect 79509 281113 79819 281147
rect 79509 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 79819 281113
rect 79509 281051 79819 281085
rect 79509 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 79819 281051
rect 79509 280989 79819 281023
rect 79509 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 79819 280989
rect 79509 272175 79819 280961
rect 79509 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 79819 272175
rect 79509 272113 79819 272147
rect 79509 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 79819 272113
rect 79509 272051 79819 272085
rect 79509 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 79819 272051
rect 79509 271989 79819 272023
rect 79509 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 79819 271989
rect 79509 263175 79819 271961
rect 79509 263147 79557 263175
rect 79585 263147 79619 263175
rect 79647 263147 79681 263175
rect 79709 263147 79743 263175
rect 79771 263147 79819 263175
rect 79509 263113 79819 263147
rect 79509 263085 79557 263113
rect 79585 263085 79619 263113
rect 79647 263085 79681 263113
rect 79709 263085 79743 263113
rect 79771 263085 79819 263113
rect 79509 263051 79819 263085
rect 79509 263023 79557 263051
rect 79585 263023 79619 263051
rect 79647 263023 79681 263051
rect 79709 263023 79743 263051
rect 79771 263023 79819 263051
rect 79509 262989 79819 263023
rect 79509 262961 79557 262989
rect 79585 262961 79619 262989
rect 79647 262961 79681 262989
rect 79709 262961 79743 262989
rect 79771 262961 79819 262989
rect 79509 254175 79819 262961
rect 79509 254147 79557 254175
rect 79585 254147 79619 254175
rect 79647 254147 79681 254175
rect 79709 254147 79743 254175
rect 79771 254147 79819 254175
rect 79509 254113 79819 254147
rect 79509 254085 79557 254113
rect 79585 254085 79619 254113
rect 79647 254085 79681 254113
rect 79709 254085 79743 254113
rect 79771 254085 79819 254113
rect 79509 254051 79819 254085
rect 79509 254023 79557 254051
rect 79585 254023 79619 254051
rect 79647 254023 79681 254051
rect 79709 254023 79743 254051
rect 79771 254023 79819 254051
rect 79509 253989 79819 254023
rect 79509 253961 79557 253989
rect 79585 253961 79619 253989
rect 79647 253961 79681 253989
rect 79709 253961 79743 253989
rect 79771 253961 79819 253989
rect 79509 245175 79819 253961
rect 79509 245147 79557 245175
rect 79585 245147 79619 245175
rect 79647 245147 79681 245175
rect 79709 245147 79743 245175
rect 79771 245147 79819 245175
rect 79509 245113 79819 245147
rect 79509 245085 79557 245113
rect 79585 245085 79619 245113
rect 79647 245085 79681 245113
rect 79709 245085 79743 245113
rect 79771 245085 79819 245113
rect 79509 245051 79819 245085
rect 79509 245023 79557 245051
rect 79585 245023 79619 245051
rect 79647 245023 79681 245051
rect 79709 245023 79743 245051
rect 79771 245023 79819 245051
rect 79509 244989 79819 245023
rect 79509 244961 79557 244989
rect 79585 244961 79619 244989
rect 79647 244961 79681 244989
rect 79709 244961 79743 244989
rect 79771 244961 79819 244989
rect 79509 236175 79819 244961
rect 79509 236147 79557 236175
rect 79585 236147 79619 236175
rect 79647 236147 79681 236175
rect 79709 236147 79743 236175
rect 79771 236147 79819 236175
rect 79509 236113 79819 236147
rect 79509 236085 79557 236113
rect 79585 236085 79619 236113
rect 79647 236085 79681 236113
rect 79709 236085 79743 236113
rect 79771 236085 79819 236113
rect 79509 236051 79819 236085
rect 79509 236023 79557 236051
rect 79585 236023 79619 236051
rect 79647 236023 79681 236051
rect 79709 236023 79743 236051
rect 79771 236023 79819 236051
rect 79509 235989 79819 236023
rect 79509 235961 79557 235989
rect 79585 235961 79619 235989
rect 79647 235961 79681 235989
rect 79709 235961 79743 235989
rect 79771 235961 79819 235989
rect 79509 227175 79819 235961
rect 79509 227147 79557 227175
rect 79585 227147 79619 227175
rect 79647 227147 79681 227175
rect 79709 227147 79743 227175
rect 79771 227147 79819 227175
rect 79509 227113 79819 227147
rect 79509 227085 79557 227113
rect 79585 227085 79619 227113
rect 79647 227085 79681 227113
rect 79709 227085 79743 227113
rect 79771 227085 79819 227113
rect 79509 227051 79819 227085
rect 79509 227023 79557 227051
rect 79585 227023 79619 227051
rect 79647 227023 79681 227051
rect 79709 227023 79743 227051
rect 79771 227023 79819 227051
rect 79509 226989 79819 227023
rect 79509 226961 79557 226989
rect 79585 226961 79619 226989
rect 79647 226961 79681 226989
rect 79709 226961 79743 226989
rect 79771 226961 79819 226989
rect 79509 218175 79819 226961
rect 79509 218147 79557 218175
rect 79585 218147 79619 218175
rect 79647 218147 79681 218175
rect 79709 218147 79743 218175
rect 79771 218147 79819 218175
rect 79509 218113 79819 218147
rect 79509 218085 79557 218113
rect 79585 218085 79619 218113
rect 79647 218085 79681 218113
rect 79709 218085 79743 218113
rect 79771 218085 79819 218113
rect 79509 218051 79819 218085
rect 79509 218023 79557 218051
rect 79585 218023 79619 218051
rect 79647 218023 79681 218051
rect 79709 218023 79743 218051
rect 79771 218023 79819 218051
rect 79509 217989 79819 218023
rect 79509 217961 79557 217989
rect 79585 217961 79619 217989
rect 79647 217961 79681 217989
rect 79709 217961 79743 217989
rect 79771 217961 79819 217989
rect 79509 209175 79819 217961
rect 79509 209147 79557 209175
rect 79585 209147 79619 209175
rect 79647 209147 79681 209175
rect 79709 209147 79743 209175
rect 79771 209147 79819 209175
rect 79509 209113 79819 209147
rect 79509 209085 79557 209113
rect 79585 209085 79619 209113
rect 79647 209085 79681 209113
rect 79709 209085 79743 209113
rect 79771 209085 79819 209113
rect 79509 209051 79819 209085
rect 79509 209023 79557 209051
rect 79585 209023 79619 209051
rect 79647 209023 79681 209051
rect 79709 209023 79743 209051
rect 79771 209023 79819 209051
rect 79509 208989 79819 209023
rect 79509 208961 79557 208989
rect 79585 208961 79619 208989
rect 79647 208961 79681 208989
rect 79709 208961 79743 208989
rect 79771 208961 79819 208989
rect 79509 200175 79819 208961
rect 79509 200147 79557 200175
rect 79585 200147 79619 200175
rect 79647 200147 79681 200175
rect 79709 200147 79743 200175
rect 79771 200147 79819 200175
rect 79509 200113 79819 200147
rect 79509 200085 79557 200113
rect 79585 200085 79619 200113
rect 79647 200085 79681 200113
rect 79709 200085 79743 200113
rect 79771 200085 79819 200113
rect 79509 200051 79819 200085
rect 79509 200023 79557 200051
rect 79585 200023 79619 200051
rect 79647 200023 79681 200051
rect 79709 200023 79743 200051
rect 79771 200023 79819 200051
rect 79509 199989 79819 200023
rect 79509 199961 79557 199989
rect 79585 199961 79619 199989
rect 79647 199961 79681 199989
rect 79709 199961 79743 199989
rect 79771 199961 79819 199989
rect 79509 191175 79819 199961
rect 79509 191147 79557 191175
rect 79585 191147 79619 191175
rect 79647 191147 79681 191175
rect 79709 191147 79743 191175
rect 79771 191147 79819 191175
rect 79509 191113 79819 191147
rect 79509 191085 79557 191113
rect 79585 191085 79619 191113
rect 79647 191085 79681 191113
rect 79709 191085 79743 191113
rect 79771 191085 79819 191113
rect 79509 191051 79819 191085
rect 79509 191023 79557 191051
rect 79585 191023 79619 191051
rect 79647 191023 79681 191051
rect 79709 191023 79743 191051
rect 79771 191023 79819 191051
rect 79509 190989 79819 191023
rect 79509 190961 79557 190989
rect 79585 190961 79619 190989
rect 79647 190961 79681 190989
rect 79709 190961 79743 190989
rect 79771 190961 79819 190989
rect 79509 182175 79819 190961
rect 79509 182147 79557 182175
rect 79585 182147 79619 182175
rect 79647 182147 79681 182175
rect 79709 182147 79743 182175
rect 79771 182147 79819 182175
rect 79509 182113 79819 182147
rect 79509 182085 79557 182113
rect 79585 182085 79619 182113
rect 79647 182085 79681 182113
rect 79709 182085 79743 182113
rect 79771 182085 79819 182113
rect 79509 182051 79819 182085
rect 79509 182023 79557 182051
rect 79585 182023 79619 182051
rect 79647 182023 79681 182051
rect 79709 182023 79743 182051
rect 79771 182023 79819 182051
rect 79509 181989 79819 182023
rect 79509 181961 79557 181989
rect 79585 181961 79619 181989
rect 79647 181961 79681 181989
rect 79709 181961 79743 181989
rect 79771 181961 79819 181989
rect 79509 173175 79819 181961
rect 79509 173147 79557 173175
rect 79585 173147 79619 173175
rect 79647 173147 79681 173175
rect 79709 173147 79743 173175
rect 79771 173147 79819 173175
rect 79509 173113 79819 173147
rect 79509 173085 79557 173113
rect 79585 173085 79619 173113
rect 79647 173085 79681 173113
rect 79709 173085 79743 173113
rect 79771 173085 79819 173113
rect 79509 173051 79819 173085
rect 79509 173023 79557 173051
rect 79585 173023 79619 173051
rect 79647 173023 79681 173051
rect 79709 173023 79743 173051
rect 79771 173023 79819 173051
rect 79509 172989 79819 173023
rect 79509 172961 79557 172989
rect 79585 172961 79619 172989
rect 79647 172961 79681 172989
rect 79709 172961 79743 172989
rect 79771 172961 79819 172989
rect 79509 164175 79819 172961
rect 79509 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 79819 164175
rect 79509 164113 79819 164147
rect 79509 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 79819 164113
rect 79509 164051 79819 164085
rect 79509 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 79819 164051
rect 79509 163989 79819 164023
rect 79509 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 79819 163989
rect 79509 155175 79819 163961
rect 79509 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 79819 155175
rect 79509 155113 79819 155147
rect 79509 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 79819 155113
rect 79509 155051 79819 155085
rect 79509 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 79819 155051
rect 79509 154989 79819 155023
rect 79509 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 79819 154989
rect 79509 146175 79819 154961
rect 79509 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 79819 146175
rect 79509 146113 79819 146147
rect 79509 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 79819 146113
rect 79509 146051 79819 146085
rect 79509 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 79819 146051
rect 79509 145989 79819 146023
rect 79509 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 79819 145989
rect 79509 137175 79819 145961
rect 79509 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 79819 137175
rect 79509 137113 79819 137147
rect 79509 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 79819 137113
rect 79509 137051 79819 137085
rect 79509 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 79819 137051
rect 79509 136989 79819 137023
rect 79509 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 79819 136989
rect 79509 128175 79819 136961
rect 79509 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 79819 128175
rect 79509 128113 79819 128147
rect 79509 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 79819 128113
rect 79509 128051 79819 128085
rect 79509 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 79819 128051
rect 79509 127989 79819 128023
rect 79509 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 79819 127989
rect 79509 119175 79819 127961
rect 79509 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 79819 119175
rect 79509 119113 79819 119147
rect 79509 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 79819 119113
rect 79509 119051 79819 119085
rect 79509 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 79819 119051
rect 79509 118989 79819 119023
rect 79509 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 79819 118989
rect 79509 110175 79819 118961
rect 79509 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 79819 110175
rect 79509 110113 79819 110147
rect 79509 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 79819 110113
rect 79509 110051 79819 110085
rect 79509 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 79819 110051
rect 79509 109989 79819 110023
rect 79509 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 79819 109989
rect 79509 101175 79819 109961
rect 79509 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 79819 101175
rect 79509 101113 79819 101147
rect 79509 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 79819 101113
rect 79509 101051 79819 101085
rect 79509 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 79819 101051
rect 79509 100989 79819 101023
rect 79509 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 79819 100989
rect 79509 92175 79819 100961
rect 79509 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 79819 92175
rect 79509 92113 79819 92147
rect 79509 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 79819 92113
rect 79509 92051 79819 92085
rect 79509 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 79819 92051
rect 79509 91989 79819 92023
rect 79509 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 79819 91989
rect 79509 83175 79819 91961
rect 79509 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 79819 83175
rect 79509 83113 79819 83147
rect 79509 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 79819 83113
rect 79509 83051 79819 83085
rect 79509 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 79819 83051
rect 79509 82989 79819 83023
rect 79509 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 79819 82989
rect 79509 74175 79819 82961
rect 79509 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 79819 74175
rect 79509 74113 79819 74147
rect 79509 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 79819 74113
rect 79509 74051 79819 74085
rect 79509 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 79819 74051
rect 79509 73989 79819 74023
rect 79509 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 79819 73989
rect 79509 65175 79819 73961
rect 79509 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 79819 65175
rect 79509 65113 79819 65147
rect 79509 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 79819 65113
rect 79509 65051 79819 65085
rect 79509 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 79819 65051
rect 79509 64989 79819 65023
rect 79509 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 79819 64989
rect 79509 56175 79819 64961
rect 79509 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 79819 56175
rect 79509 56113 79819 56147
rect 79509 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 79819 56113
rect 79509 56051 79819 56085
rect 79509 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 79819 56051
rect 79509 55989 79819 56023
rect 79509 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 79819 55989
rect 79509 47175 79819 55961
rect 79509 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 79819 47175
rect 79509 47113 79819 47147
rect 79509 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 79819 47113
rect 79509 47051 79819 47085
rect 79509 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 79819 47051
rect 79509 46989 79819 47023
rect 79509 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 79819 46989
rect 79509 38175 79819 46961
rect 79509 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 79819 38175
rect 79509 38113 79819 38147
rect 79509 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 79819 38113
rect 79509 38051 79819 38085
rect 79509 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 79819 38051
rect 79509 37989 79819 38023
rect 79509 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 79819 37989
rect 79509 29175 79819 37961
rect 79509 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 79819 29175
rect 79509 29113 79819 29147
rect 79509 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 79819 29113
rect 79509 29051 79819 29085
rect 79509 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 79819 29051
rect 79509 28989 79819 29023
rect 79509 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 79819 28989
rect 79509 20175 79819 28961
rect 79509 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 79819 20175
rect 79509 20113 79819 20147
rect 79509 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 79819 20113
rect 79509 20051 79819 20085
rect 79509 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 79819 20051
rect 79509 19989 79819 20023
rect 79509 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 79819 19989
rect 79509 11175 79819 19961
rect 79509 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 79819 11175
rect 79509 11113 79819 11147
rect 79509 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 79819 11113
rect 79509 11051 79819 11085
rect 79509 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 79819 11051
rect 79509 10989 79819 11023
rect 79509 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 79819 10989
rect 79509 2175 79819 10961
rect 79509 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 79819 2175
rect 79509 2113 79819 2147
rect 79509 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 79819 2113
rect 79509 2051 79819 2085
rect 79509 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 79819 2051
rect 79509 1989 79819 2023
rect 79509 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 79819 1989
rect 79509 -80 79819 1961
rect 79509 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 79819 -80
rect 79509 -142 79819 -108
rect 79509 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 79819 -142
rect 79509 -204 79819 -170
rect 79509 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 79819 -204
rect 79509 -266 79819 -232
rect 79509 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 79819 -266
rect 79509 -822 79819 -294
rect 81369 299086 81679 299134
rect 81369 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 81679 299086
rect 81369 299024 81679 299058
rect 81369 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 81679 299024
rect 81369 298962 81679 298996
rect 81369 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 81679 298962
rect 81369 298900 81679 298934
rect 81369 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 81679 298900
rect 81369 293175 81679 298872
rect 81369 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 81679 293175
rect 81369 293113 81679 293147
rect 81369 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 81679 293113
rect 81369 293051 81679 293085
rect 81369 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 81679 293051
rect 81369 292989 81679 293023
rect 81369 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 81679 292989
rect 81369 284175 81679 292961
rect 81369 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 81679 284175
rect 81369 284113 81679 284147
rect 81369 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 81679 284113
rect 81369 284051 81679 284085
rect 81369 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 81679 284051
rect 81369 283989 81679 284023
rect 81369 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 81679 283989
rect 81369 275175 81679 283961
rect 81369 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 81679 275175
rect 81369 275113 81679 275147
rect 81369 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 81679 275113
rect 81369 275051 81679 275085
rect 81369 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 81679 275051
rect 81369 274989 81679 275023
rect 81369 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 81679 274989
rect 81369 266175 81679 274961
rect 81369 266147 81417 266175
rect 81445 266147 81479 266175
rect 81507 266147 81541 266175
rect 81569 266147 81603 266175
rect 81631 266147 81679 266175
rect 81369 266113 81679 266147
rect 81369 266085 81417 266113
rect 81445 266085 81479 266113
rect 81507 266085 81541 266113
rect 81569 266085 81603 266113
rect 81631 266085 81679 266113
rect 81369 266051 81679 266085
rect 81369 266023 81417 266051
rect 81445 266023 81479 266051
rect 81507 266023 81541 266051
rect 81569 266023 81603 266051
rect 81631 266023 81679 266051
rect 81369 265989 81679 266023
rect 81369 265961 81417 265989
rect 81445 265961 81479 265989
rect 81507 265961 81541 265989
rect 81569 265961 81603 265989
rect 81631 265961 81679 265989
rect 81369 257175 81679 265961
rect 81369 257147 81417 257175
rect 81445 257147 81479 257175
rect 81507 257147 81541 257175
rect 81569 257147 81603 257175
rect 81631 257147 81679 257175
rect 81369 257113 81679 257147
rect 81369 257085 81417 257113
rect 81445 257085 81479 257113
rect 81507 257085 81541 257113
rect 81569 257085 81603 257113
rect 81631 257085 81679 257113
rect 81369 257051 81679 257085
rect 81369 257023 81417 257051
rect 81445 257023 81479 257051
rect 81507 257023 81541 257051
rect 81569 257023 81603 257051
rect 81631 257023 81679 257051
rect 81369 256989 81679 257023
rect 81369 256961 81417 256989
rect 81445 256961 81479 256989
rect 81507 256961 81541 256989
rect 81569 256961 81603 256989
rect 81631 256961 81679 256989
rect 81369 248175 81679 256961
rect 81369 248147 81417 248175
rect 81445 248147 81479 248175
rect 81507 248147 81541 248175
rect 81569 248147 81603 248175
rect 81631 248147 81679 248175
rect 81369 248113 81679 248147
rect 81369 248085 81417 248113
rect 81445 248085 81479 248113
rect 81507 248085 81541 248113
rect 81569 248085 81603 248113
rect 81631 248085 81679 248113
rect 81369 248051 81679 248085
rect 81369 248023 81417 248051
rect 81445 248023 81479 248051
rect 81507 248023 81541 248051
rect 81569 248023 81603 248051
rect 81631 248023 81679 248051
rect 81369 247989 81679 248023
rect 81369 247961 81417 247989
rect 81445 247961 81479 247989
rect 81507 247961 81541 247989
rect 81569 247961 81603 247989
rect 81631 247961 81679 247989
rect 81369 239175 81679 247961
rect 81369 239147 81417 239175
rect 81445 239147 81479 239175
rect 81507 239147 81541 239175
rect 81569 239147 81603 239175
rect 81631 239147 81679 239175
rect 81369 239113 81679 239147
rect 81369 239085 81417 239113
rect 81445 239085 81479 239113
rect 81507 239085 81541 239113
rect 81569 239085 81603 239113
rect 81631 239085 81679 239113
rect 81369 239051 81679 239085
rect 81369 239023 81417 239051
rect 81445 239023 81479 239051
rect 81507 239023 81541 239051
rect 81569 239023 81603 239051
rect 81631 239023 81679 239051
rect 81369 238989 81679 239023
rect 81369 238961 81417 238989
rect 81445 238961 81479 238989
rect 81507 238961 81541 238989
rect 81569 238961 81603 238989
rect 81631 238961 81679 238989
rect 81369 230175 81679 238961
rect 81369 230147 81417 230175
rect 81445 230147 81479 230175
rect 81507 230147 81541 230175
rect 81569 230147 81603 230175
rect 81631 230147 81679 230175
rect 81369 230113 81679 230147
rect 81369 230085 81417 230113
rect 81445 230085 81479 230113
rect 81507 230085 81541 230113
rect 81569 230085 81603 230113
rect 81631 230085 81679 230113
rect 81369 230051 81679 230085
rect 81369 230023 81417 230051
rect 81445 230023 81479 230051
rect 81507 230023 81541 230051
rect 81569 230023 81603 230051
rect 81631 230023 81679 230051
rect 81369 229989 81679 230023
rect 81369 229961 81417 229989
rect 81445 229961 81479 229989
rect 81507 229961 81541 229989
rect 81569 229961 81603 229989
rect 81631 229961 81679 229989
rect 81369 221175 81679 229961
rect 81369 221147 81417 221175
rect 81445 221147 81479 221175
rect 81507 221147 81541 221175
rect 81569 221147 81603 221175
rect 81631 221147 81679 221175
rect 81369 221113 81679 221147
rect 81369 221085 81417 221113
rect 81445 221085 81479 221113
rect 81507 221085 81541 221113
rect 81569 221085 81603 221113
rect 81631 221085 81679 221113
rect 81369 221051 81679 221085
rect 81369 221023 81417 221051
rect 81445 221023 81479 221051
rect 81507 221023 81541 221051
rect 81569 221023 81603 221051
rect 81631 221023 81679 221051
rect 81369 220989 81679 221023
rect 81369 220961 81417 220989
rect 81445 220961 81479 220989
rect 81507 220961 81541 220989
rect 81569 220961 81603 220989
rect 81631 220961 81679 220989
rect 81369 212175 81679 220961
rect 81369 212147 81417 212175
rect 81445 212147 81479 212175
rect 81507 212147 81541 212175
rect 81569 212147 81603 212175
rect 81631 212147 81679 212175
rect 81369 212113 81679 212147
rect 81369 212085 81417 212113
rect 81445 212085 81479 212113
rect 81507 212085 81541 212113
rect 81569 212085 81603 212113
rect 81631 212085 81679 212113
rect 81369 212051 81679 212085
rect 81369 212023 81417 212051
rect 81445 212023 81479 212051
rect 81507 212023 81541 212051
rect 81569 212023 81603 212051
rect 81631 212023 81679 212051
rect 81369 211989 81679 212023
rect 81369 211961 81417 211989
rect 81445 211961 81479 211989
rect 81507 211961 81541 211989
rect 81569 211961 81603 211989
rect 81631 211961 81679 211989
rect 81369 203175 81679 211961
rect 81369 203147 81417 203175
rect 81445 203147 81479 203175
rect 81507 203147 81541 203175
rect 81569 203147 81603 203175
rect 81631 203147 81679 203175
rect 81369 203113 81679 203147
rect 81369 203085 81417 203113
rect 81445 203085 81479 203113
rect 81507 203085 81541 203113
rect 81569 203085 81603 203113
rect 81631 203085 81679 203113
rect 81369 203051 81679 203085
rect 81369 203023 81417 203051
rect 81445 203023 81479 203051
rect 81507 203023 81541 203051
rect 81569 203023 81603 203051
rect 81631 203023 81679 203051
rect 81369 202989 81679 203023
rect 81369 202961 81417 202989
rect 81445 202961 81479 202989
rect 81507 202961 81541 202989
rect 81569 202961 81603 202989
rect 81631 202961 81679 202989
rect 81369 194175 81679 202961
rect 81369 194147 81417 194175
rect 81445 194147 81479 194175
rect 81507 194147 81541 194175
rect 81569 194147 81603 194175
rect 81631 194147 81679 194175
rect 81369 194113 81679 194147
rect 81369 194085 81417 194113
rect 81445 194085 81479 194113
rect 81507 194085 81541 194113
rect 81569 194085 81603 194113
rect 81631 194085 81679 194113
rect 81369 194051 81679 194085
rect 81369 194023 81417 194051
rect 81445 194023 81479 194051
rect 81507 194023 81541 194051
rect 81569 194023 81603 194051
rect 81631 194023 81679 194051
rect 81369 193989 81679 194023
rect 81369 193961 81417 193989
rect 81445 193961 81479 193989
rect 81507 193961 81541 193989
rect 81569 193961 81603 193989
rect 81631 193961 81679 193989
rect 81369 185175 81679 193961
rect 81369 185147 81417 185175
rect 81445 185147 81479 185175
rect 81507 185147 81541 185175
rect 81569 185147 81603 185175
rect 81631 185147 81679 185175
rect 81369 185113 81679 185147
rect 81369 185085 81417 185113
rect 81445 185085 81479 185113
rect 81507 185085 81541 185113
rect 81569 185085 81603 185113
rect 81631 185085 81679 185113
rect 81369 185051 81679 185085
rect 81369 185023 81417 185051
rect 81445 185023 81479 185051
rect 81507 185023 81541 185051
rect 81569 185023 81603 185051
rect 81631 185023 81679 185051
rect 81369 184989 81679 185023
rect 81369 184961 81417 184989
rect 81445 184961 81479 184989
rect 81507 184961 81541 184989
rect 81569 184961 81603 184989
rect 81631 184961 81679 184989
rect 81369 176175 81679 184961
rect 81369 176147 81417 176175
rect 81445 176147 81479 176175
rect 81507 176147 81541 176175
rect 81569 176147 81603 176175
rect 81631 176147 81679 176175
rect 81369 176113 81679 176147
rect 81369 176085 81417 176113
rect 81445 176085 81479 176113
rect 81507 176085 81541 176113
rect 81569 176085 81603 176113
rect 81631 176085 81679 176113
rect 81369 176051 81679 176085
rect 81369 176023 81417 176051
rect 81445 176023 81479 176051
rect 81507 176023 81541 176051
rect 81569 176023 81603 176051
rect 81631 176023 81679 176051
rect 81369 175989 81679 176023
rect 81369 175961 81417 175989
rect 81445 175961 81479 175989
rect 81507 175961 81541 175989
rect 81569 175961 81603 175989
rect 81631 175961 81679 175989
rect 81369 167175 81679 175961
rect 81369 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 81679 167175
rect 81369 167113 81679 167147
rect 81369 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 81679 167113
rect 81369 167051 81679 167085
rect 81369 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 81679 167051
rect 81369 166989 81679 167023
rect 81369 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 81679 166989
rect 81369 158175 81679 166961
rect 81369 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 81679 158175
rect 81369 158113 81679 158147
rect 81369 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 81679 158113
rect 81369 158051 81679 158085
rect 81369 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 81679 158051
rect 81369 157989 81679 158023
rect 81369 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 81679 157989
rect 81369 149175 81679 157961
rect 81369 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 81679 149175
rect 81369 149113 81679 149147
rect 81369 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 81679 149113
rect 81369 149051 81679 149085
rect 81369 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 81679 149051
rect 81369 148989 81679 149023
rect 81369 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 81679 148989
rect 81369 140175 81679 148961
rect 81369 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 81679 140175
rect 81369 140113 81679 140147
rect 81369 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 81679 140113
rect 81369 140051 81679 140085
rect 81369 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 81679 140051
rect 81369 139989 81679 140023
rect 81369 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 81679 139989
rect 81369 131175 81679 139961
rect 81369 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 81679 131175
rect 81369 131113 81679 131147
rect 81369 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 81679 131113
rect 81369 131051 81679 131085
rect 81369 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 81679 131051
rect 81369 130989 81679 131023
rect 81369 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 81679 130989
rect 81369 122175 81679 130961
rect 81369 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 81679 122175
rect 81369 122113 81679 122147
rect 81369 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 81679 122113
rect 81369 122051 81679 122085
rect 81369 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 81679 122051
rect 81369 121989 81679 122023
rect 81369 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 81679 121989
rect 81369 113175 81679 121961
rect 81369 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 81679 113175
rect 81369 113113 81679 113147
rect 81369 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 81679 113113
rect 81369 113051 81679 113085
rect 81369 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 81679 113051
rect 81369 112989 81679 113023
rect 81369 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 81679 112989
rect 81369 104175 81679 112961
rect 81369 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 81679 104175
rect 81369 104113 81679 104147
rect 81369 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 81679 104113
rect 81369 104051 81679 104085
rect 81369 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 81679 104051
rect 81369 103989 81679 104023
rect 81369 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 81679 103989
rect 81369 95175 81679 103961
rect 81369 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 81679 95175
rect 81369 95113 81679 95147
rect 81369 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 81679 95113
rect 81369 95051 81679 95085
rect 81369 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 81679 95051
rect 81369 94989 81679 95023
rect 81369 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 81679 94989
rect 81369 86175 81679 94961
rect 81369 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 81679 86175
rect 81369 86113 81679 86147
rect 81369 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 81679 86113
rect 81369 86051 81679 86085
rect 81369 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 81679 86051
rect 81369 85989 81679 86023
rect 81369 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 81679 85989
rect 81369 77175 81679 85961
rect 81369 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 81679 77175
rect 81369 77113 81679 77147
rect 81369 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 81679 77113
rect 81369 77051 81679 77085
rect 81369 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 81679 77051
rect 81369 76989 81679 77023
rect 81369 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 81679 76989
rect 81369 68175 81679 76961
rect 81369 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 81679 68175
rect 81369 68113 81679 68147
rect 81369 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 81679 68113
rect 81369 68051 81679 68085
rect 81369 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 81679 68051
rect 81369 67989 81679 68023
rect 81369 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 81679 67989
rect 81369 59175 81679 67961
rect 81369 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 81679 59175
rect 81369 59113 81679 59147
rect 81369 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 81679 59113
rect 81369 59051 81679 59085
rect 81369 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 81679 59051
rect 81369 58989 81679 59023
rect 81369 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 81679 58989
rect 81369 50175 81679 58961
rect 81369 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 81679 50175
rect 81369 50113 81679 50147
rect 81369 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 81679 50113
rect 81369 50051 81679 50085
rect 81369 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 81679 50051
rect 81369 49989 81679 50023
rect 81369 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 81679 49989
rect 81369 41175 81679 49961
rect 81369 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 81679 41175
rect 81369 41113 81679 41147
rect 81369 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 81679 41113
rect 81369 41051 81679 41085
rect 81369 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 81679 41051
rect 81369 40989 81679 41023
rect 81369 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 81679 40989
rect 81369 32175 81679 40961
rect 81369 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 81679 32175
rect 81369 32113 81679 32147
rect 81369 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 81679 32113
rect 81369 32051 81679 32085
rect 81369 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 81679 32051
rect 81369 31989 81679 32023
rect 81369 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 81679 31989
rect 81369 23175 81679 31961
rect 81369 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 81679 23175
rect 81369 23113 81679 23147
rect 81369 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 81679 23113
rect 81369 23051 81679 23085
rect 81369 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 81679 23051
rect 81369 22989 81679 23023
rect 81369 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 81679 22989
rect 81369 14175 81679 22961
rect 81369 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 81679 14175
rect 81369 14113 81679 14147
rect 81369 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 81679 14113
rect 81369 14051 81679 14085
rect 81369 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 81679 14051
rect 81369 13989 81679 14023
rect 81369 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 81679 13989
rect 81369 5175 81679 13961
rect 81369 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 81679 5175
rect 81369 5113 81679 5147
rect 81369 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 81679 5113
rect 81369 5051 81679 5085
rect 81369 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 81679 5051
rect 81369 4989 81679 5023
rect 81369 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 81679 4989
rect 81369 -560 81679 4961
rect 81369 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 81679 -560
rect 81369 -622 81679 -588
rect 81369 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 81679 -622
rect 81369 -684 81679 -650
rect 81369 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 81679 -684
rect 81369 -746 81679 -712
rect 81369 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 81679 -746
rect 81369 -822 81679 -774
rect 94869 298606 95179 299134
rect 94869 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 95179 298606
rect 94869 298544 95179 298578
rect 94869 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 95179 298544
rect 94869 298482 95179 298516
rect 94869 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 95179 298482
rect 94869 298420 95179 298454
rect 94869 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 95179 298420
rect 94869 290175 95179 298392
rect 94869 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 95179 290175
rect 94869 290113 95179 290147
rect 94869 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 95179 290113
rect 94869 290051 95179 290085
rect 94869 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 95179 290051
rect 94869 289989 95179 290023
rect 94869 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 95179 289989
rect 94869 281175 95179 289961
rect 94869 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 95179 281175
rect 94869 281113 95179 281147
rect 94869 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 95179 281113
rect 94869 281051 95179 281085
rect 94869 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 95179 281051
rect 94869 280989 95179 281023
rect 94869 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 95179 280989
rect 94869 272175 95179 280961
rect 94869 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 95179 272175
rect 94869 272113 95179 272147
rect 94869 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 95179 272113
rect 94869 272051 95179 272085
rect 94869 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 95179 272051
rect 94869 271989 95179 272023
rect 94869 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 95179 271989
rect 94869 263175 95179 271961
rect 94869 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 95179 263175
rect 94869 263113 95179 263147
rect 94869 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 95179 263113
rect 94869 263051 95179 263085
rect 94869 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 95179 263051
rect 94869 262989 95179 263023
rect 94869 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 95179 262989
rect 94869 254175 95179 262961
rect 94869 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 95179 254175
rect 94869 254113 95179 254147
rect 94869 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 95179 254113
rect 94869 254051 95179 254085
rect 94869 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 95179 254051
rect 94869 253989 95179 254023
rect 94869 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 95179 253989
rect 94869 245175 95179 253961
rect 94869 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 95179 245175
rect 94869 245113 95179 245147
rect 94869 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 95179 245113
rect 94869 245051 95179 245085
rect 94869 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 95179 245051
rect 94869 244989 95179 245023
rect 94869 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 95179 244989
rect 94869 236175 95179 244961
rect 94869 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 95179 236175
rect 94869 236113 95179 236147
rect 94869 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 95179 236113
rect 94869 236051 95179 236085
rect 94869 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 95179 236051
rect 94869 235989 95179 236023
rect 94869 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 95179 235989
rect 94869 227175 95179 235961
rect 94869 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 95179 227175
rect 94869 227113 95179 227147
rect 94869 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 95179 227113
rect 94869 227051 95179 227085
rect 94869 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 95179 227051
rect 94869 226989 95179 227023
rect 94869 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 95179 226989
rect 94869 218175 95179 226961
rect 94869 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 95179 218175
rect 94869 218113 95179 218147
rect 94869 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 95179 218113
rect 94869 218051 95179 218085
rect 94869 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 95179 218051
rect 94869 217989 95179 218023
rect 94869 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 95179 217989
rect 94869 209175 95179 217961
rect 94869 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 95179 209175
rect 94869 209113 95179 209147
rect 94869 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 95179 209113
rect 94869 209051 95179 209085
rect 94869 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 95179 209051
rect 94869 208989 95179 209023
rect 94869 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 95179 208989
rect 94869 200175 95179 208961
rect 94869 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 95179 200175
rect 94869 200113 95179 200147
rect 94869 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 95179 200113
rect 94869 200051 95179 200085
rect 94869 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 95179 200051
rect 94869 199989 95179 200023
rect 94869 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 95179 199989
rect 94869 191175 95179 199961
rect 94869 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 95179 191175
rect 94869 191113 95179 191147
rect 94869 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 95179 191113
rect 94869 191051 95179 191085
rect 94869 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 95179 191051
rect 94869 190989 95179 191023
rect 94869 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 95179 190989
rect 94869 182175 95179 190961
rect 94869 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 95179 182175
rect 94869 182113 95179 182147
rect 94869 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 95179 182113
rect 94869 182051 95179 182085
rect 94869 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 95179 182051
rect 94869 181989 95179 182023
rect 94869 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 95179 181989
rect 94869 173175 95179 181961
rect 94869 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 95179 173175
rect 94869 173113 95179 173147
rect 94869 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 95179 173113
rect 94869 173051 95179 173085
rect 94869 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 95179 173051
rect 94869 172989 95179 173023
rect 94869 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 95179 172989
rect 94869 164175 95179 172961
rect 94869 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 95179 164175
rect 94869 164113 95179 164147
rect 94869 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 95179 164113
rect 94869 164051 95179 164085
rect 94869 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 95179 164051
rect 94869 163989 95179 164023
rect 94869 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 95179 163989
rect 94869 155175 95179 163961
rect 94869 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 95179 155175
rect 94869 155113 95179 155147
rect 94869 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 95179 155113
rect 94869 155051 95179 155085
rect 94869 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 95179 155051
rect 94869 154989 95179 155023
rect 94869 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 95179 154989
rect 94869 146175 95179 154961
rect 94869 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 95179 146175
rect 94869 146113 95179 146147
rect 94869 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 95179 146113
rect 94869 146051 95179 146085
rect 94869 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 95179 146051
rect 94869 145989 95179 146023
rect 94869 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 95179 145989
rect 94869 137175 95179 145961
rect 94869 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 95179 137175
rect 94869 137113 95179 137147
rect 94869 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 95179 137113
rect 94869 137051 95179 137085
rect 94869 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 95179 137051
rect 94869 136989 95179 137023
rect 94869 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 95179 136989
rect 94869 128175 95179 136961
rect 94869 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 95179 128175
rect 94869 128113 95179 128147
rect 94869 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 95179 128113
rect 94869 128051 95179 128085
rect 94869 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 95179 128051
rect 94869 127989 95179 128023
rect 94869 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 95179 127989
rect 94869 119175 95179 127961
rect 94869 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 95179 119175
rect 94869 119113 95179 119147
rect 94869 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 95179 119113
rect 94869 119051 95179 119085
rect 94869 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 95179 119051
rect 94869 118989 95179 119023
rect 94869 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 95179 118989
rect 94869 110175 95179 118961
rect 94869 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 95179 110175
rect 94869 110113 95179 110147
rect 94869 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 95179 110113
rect 94869 110051 95179 110085
rect 94869 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 95179 110051
rect 94869 109989 95179 110023
rect 94869 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 95179 109989
rect 94869 101175 95179 109961
rect 94869 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 95179 101175
rect 94869 101113 95179 101147
rect 94869 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 95179 101113
rect 94869 101051 95179 101085
rect 94869 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 95179 101051
rect 94869 100989 95179 101023
rect 94869 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 95179 100989
rect 94869 92175 95179 100961
rect 94869 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 95179 92175
rect 94869 92113 95179 92147
rect 94869 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 95179 92113
rect 94869 92051 95179 92085
rect 94869 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 95179 92051
rect 94869 91989 95179 92023
rect 94869 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 95179 91989
rect 94869 83175 95179 91961
rect 94869 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 95179 83175
rect 94869 83113 95179 83147
rect 94869 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 95179 83113
rect 94869 83051 95179 83085
rect 94869 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 95179 83051
rect 94869 82989 95179 83023
rect 94869 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 95179 82989
rect 94869 74175 95179 82961
rect 94869 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 95179 74175
rect 94869 74113 95179 74147
rect 94869 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 95179 74113
rect 94869 74051 95179 74085
rect 94869 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 95179 74051
rect 94869 73989 95179 74023
rect 94869 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 95179 73989
rect 94869 65175 95179 73961
rect 94869 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 95179 65175
rect 94869 65113 95179 65147
rect 94869 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 95179 65113
rect 94869 65051 95179 65085
rect 94869 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 95179 65051
rect 94869 64989 95179 65023
rect 94869 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 95179 64989
rect 94869 56175 95179 64961
rect 94869 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 95179 56175
rect 94869 56113 95179 56147
rect 94869 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 95179 56113
rect 94869 56051 95179 56085
rect 94869 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 95179 56051
rect 94869 55989 95179 56023
rect 94869 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 95179 55989
rect 94869 47175 95179 55961
rect 94869 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 95179 47175
rect 94869 47113 95179 47147
rect 94869 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 95179 47113
rect 94869 47051 95179 47085
rect 94869 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 95179 47051
rect 94869 46989 95179 47023
rect 94869 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 95179 46989
rect 94869 38175 95179 46961
rect 94869 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 95179 38175
rect 94869 38113 95179 38147
rect 94869 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 95179 38113
rect 94869 38051 95179 38085
rect 94869 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 95179 38051
rect 94869 37989 95179 38023
rect 94869 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 95179 37989
rect 94869 29175 95179 37961
rect 94869 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 95179 29175
rect 94869 29113 95179 29147
rect 94869 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 95179 29113
rect 94869 29051 95179 29085
rect 94869 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 95179 29051
rect 94869 28989 95179 29023
rect 94869 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 95179 28989
rect 94869 20175 95179 28961
rect 94869 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 95179 20175
rect 94869 20113 95179 20147
rect 94869 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 95179 20113
rect 94869 20051 95179 20085
rect 94869 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 95179 20051
rect 94869 19989 95179 20023
rect 94869 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 95179 19989
rect 94869 11175 95179 19961
rect 94869 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 95179 11175
rect 94869 11113 95179 11147
rect 94869 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 95179 11113
rect 94869 11051 95179 11085
rect 94869 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 95179 11051
rect 94869 10989 95179 11023
rect 94869 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 95179 10989
rect 94869 2175 95179 10961
rect 94869 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 95179 2175
rect 94869 2113 95179 2147
rect 94869 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 95179 2113
rect 94869 2051 95179 2085
rect 94869 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 95179 2051
rect 94869 1989 95179 2023
rect 94869 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 95179 1989
rect 94869 -80 95179 1961
rect 94869 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 95179 -80
rect 94869 -142 95179 -108
rect 94869 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 95179 -142
rect 94869 -204 95179 -170
rect 94869 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 95179 -204
rect 94869 -266 95179 -232
rect 94869 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 95179 -266
rect 94869 -822 95179 -294
rect 96729 299086 97039 299134
rect 96729 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 97039 299086
rect 96729 299024 97039 299058
rect 96729 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 97039 299024
rect 96729 298962 97039 298996
rect 96729 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 97039 298962
rect 96729 298900 97039 298934
rect 96729 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 97039 298900
rect 96729 293175 97039 298872
rect 96729 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 97039 293175
rect 96729 293113 97039 293147
rect 96729 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 97039 293113
rect 96729 293051 97039 293085
rect 96729 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 97039 293051
rect 96729 292989 97039 293023
rect 96729 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 97039 292989
rect 96729 284175 97039 292961
rect 96729 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 97039 284175
rect 96729 284113 97039 284147
rect 96729 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 97039 284113
rect 96729 284051 97039 284085
rect 96729 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 97039 284051
rect 96729 283989 97039 284023
rect 96729 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 97039 283989
rect 96729 275175 97039 283961
rect 110229 298606 110539 299134
rect 110229 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 110539 298606
rect 110229 298544 110539 298578
rect 110229 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 110539 298544
rect 110229 298482 110539 298516
rect 110229 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 110539 298482
rect 110229 298420 110539 298454
rect 110229 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 110539 298420
rect 110229 290175 110539 298392
rect 110229 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 110539 290175
rect 110229 290113 110539 290147
rect 110229 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 110539 290113
rect 110229 290051 110539 290085
rect 110229 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 110539 290051
rect 110229 289989 110539 290023
rect 110229 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 110539 289989
rect 110229 281175 110539 289961
rect 110229 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 110539 281175
rect 110229 281113 110539 281147
rect 110229 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 110539 281113
rect 110229 281051 110539 281085
rect 110229 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 110539 281051
rect 110229 280989 110539 281023
rect 110229 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 110539 280989
rect 110229 276831 110539 280961
rect 112089 299086 112399 299134
rect 112089 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 112399 299086
rect 112089 299024 112399 299058
rect 112089 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 112399 299024
rect 112089 298962 112399 298996
rect 112089 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 112399 298962
rect 112089 298900 112399 298934
rect 112089 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 112399 298900
rect 112089 293175 112399 298872
rect 112089 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 112399 293175
rect 112089 293113 112399 293147
rect 112089 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 112399 293113
rect 112089 293051 112399 293085
rect 112089 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 112399 293051
rect 112089 292989 112399 293023
rect 112089 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 112399 292989
rect 112089 284175 112399 292961
rect 112089 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 112399 284175
rect 112089 284113 112399 284147
rect 112089 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 112399 284113
rect 112089 284051 112399 284085
rect 112089 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 112399 284051
rect 112089 283989 112399 284023
rect 112089 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 112399 283989
rect 112089 276831 112399 283961
rect 125589 298606 125899 299134
rect 125589 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 125899 298606
rect 125589 298544 125899 298578
rect 125589 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 125899 298544
rect 125589 298482 125899 298516
rect 125589 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 125899 298482
rect 125589 298420 125899 298454
rect 125589 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 125899 298420
rect 125589 290175 125899 298392
rect 125589 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 125899 290175
rect 125589 290113 125899 290147
rect 125589 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 125899 290113
rect 125589 290051 125899 290085
rect 125589 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 125899 290051
rect 125589 289989 125899 290023
rect 125589 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 125899 289989
rect 125589 281175 125899 289961
rect 125589 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 125899 281175
rect 125589 281113 125899 281147
rect 125589 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 125899 281113
rect 125589 281051 125899 281085
rect 125589 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 125899 281051
rect 125589 280989 125899 281023
rect 125589 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 125899 280989
rect 125589 276831 125899 280961
rect 127449 299086 127759 299134
rect 127449 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 127759 299086
rect 127449 299024 127759 299058
rect 127449 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 127759 299024
rect 127449 298962 127759 298996
rect 127449 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 127759 298962
rect 127449 298900 127759 298934
rect 127449 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 127759 298900
rect 127449 293175 127759 298872
rect 127449 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 127759 293175
rect 127449 293113 127759 293147
rect 127449 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 127759 293113
rect 127449 293051 127759 293085
rect 127449 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 127759 293051
rect 127449 292989 127759 293023
rect 127449 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 127759 292989
rect 127449 284175 127759 292961
rect 127449 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 127759 284175
rect 127449 284113 127759 284147
rect 127449 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 127759 284113
rect 127449 284051 127759 284085
rect 127449 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 127759 284051
rect 127449 283989 127759 284023
rect 127449 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 127759 283989
rect 127449 276831 127759 283961
rect 140949 298606 141259 299134
rect 140949 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 141259 298606
rect 140949 298544 141259 298578
rect 140949 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 141259 298544
rect 140949 298482 141259 298516
rect 140949 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 141259 298482
rect 140949 298420 141259 298454
rect 140949 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 141259 298420
rect 140949 290175 141259 298392
rect 140949 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 141259 290175
rect 140949 290113 141259 290147
rect 140949 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 141259 290113
rect 140949 290051 141259 290085
rect 140949 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 141259 290051
rect 140949 289989 141259 290023
rect 140949 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 141259 289989
rect 140949 281175 141259 289961
rect 140949 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 141259 281175
rect 140949 281113 141259 281147
rect 140949 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 141259 281113
rect 140949 281051 141259 281085
rect 140949 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 141259 281051
rect 140949 280989 141259 281023
rect 140949 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 141259 280989
rect 140949 276831 141259 280961
rect 142809 299086 143119 299134
rect 142809 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 143119 299086
rect 142809 299024 143119 299058
rect 142809 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 143119 299024
rect 142809 298962 143119 298996
rect 142809 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 143119 298962
rect 142809 298900 143119 298934
rect 142809 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 143119 298900
rect 142809 293175 143119 298872
rect 142809 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 143119 293175
rect 142809 293113 143119 293147
rect 142809 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 143119 293113
rect 142809 293051 143119 293085
rect 142809 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 143119 293051
rect 142809 292989 143119 293023
rect 142809 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 143119 292989
rect 142809 284175 143119 292961
rect 142809 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 143119 284175
rect 142809 284113 143119 284147
rect 142809 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 143119 284113
rect 142809 284051 143119 284085
rect 142809 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 143119 284051
rect 142809 283989 143119 284023
rect 142809 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 143119 283989
rect 142809 276831 143119 283961
rect 156309 298606 156619 299134
rect 156309 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 156619 298606
rect 156309 298544 156619 298578
rect 156309 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 156619 298544
rect 156309 298482 156619 298516
rect 156309 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 156619 298482
rect 156309 298420 156619 298454
rect 156309 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 156619 298420
rect 156309 290175 156619 298392
rect 156309 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 156619 290175
rect 156309 290113 156619 290147
rect 156309 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 156619 290113
rect 156309 290051 156619 290085
rect 156309 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 156619 290051
rect 156309 289989 156619 290023
rect 156309 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 156619 289989
rect 156309 281175 156619 289961
rect 156309 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 156619 281175
rect 156309 281113 156619 281147
rect 156309 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 156619 281113
rect 156309 281051 156619 281085
rect 156309 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 156619 281051
rect 156309 280989 156619 281023
rect 156309 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 156619 280989
rect 156309 276831 156619 280961
rect 158169 299086 158479 299134
rect 158169 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 158479 299086
rect 158169 299024 158479 299058
rect 158169 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 158479 299024
rect 158169 298962 158479 298996
rect 158169 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 158479 298962
rect 158169 298900 158479 298934
rect 158169 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 158479 298900
rect 158169 293175 158479 298872
rect 158169 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 158479 293175
rect 158169 293113 158479 293147
rect 158169 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 158479 293113
rect 158169 293051 158479 293085
rect 158169 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 158479 293051
rect 158169 292989 158479 293023
rect 158169 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 158479 292989
rect 158169 284175 158479 292961
rect 158169 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 158479 284175
rect 158169 284113 158479 284147
rect 158169 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 158479 284113
rect 158169 284051 158479 284085
rect 158169 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 158479 284051
rect 158169 283989 158479 284023
rect 158169 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 158479 283989
rect 158169 276831 158479 283961
rect 171669 298606 171979 299134
rect 171669 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 171979 298606
rect 171669 298544 171979 298578
rect 171669 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 171979 298544
rect 171669 298482 171979 298516
rect 171669 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 171979 298482
rect 171669 298420 171979 298454
rect 171669 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 171979 298420
rect 171669 290175 171979 298392
rect 171669 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 171979 290175
rect 171669 290113 171979 290147
rect 171669 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 171979 290113
rect 171669 290051 171979 290085
rect 171669 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 171979 290051
rect 171669 289989 171979 290023
rect 171669 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 171979 289989
rect 171669 281175 171979 289961
rect 171669 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 171979 281175
rect 171669 281113 171979 281147
rect 171669 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 171979 281113
rect 171669 281051 171979 281085
rect 171669 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 171979 281051
rect 171669 280989 171979 281023
rect 171669 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 171979 280989
rect 171669 276831 171979 280961
rect 173529 299086 173839 299134
rect 173529 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 173839 299086
rect 173529 299024 173839 299058
rect 173529 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 173839 299024
rect 173529 298962 173839 298996
rect 173529 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 173839 298962
rect 173529 298900 173839 298934
rect 173529 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 173839 298900
rect 173529 293175 173839 298872
rect 173529 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 173839 293175
rect 173529 293113 173839 293147
rect 173529 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 173839 293113
rect 173529 293051 173839 293085
rect 173529 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 173839 293051
rect 173529 292989 173839 293023
rect 173529 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 173839 292989
rect 173529 284175 173839 292961
rect 173529 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 173839 284175
rect 173529 284113 173839 284147
rect 173529 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 173839 284113
rect 173529 284051 173839 284085
rect 173529 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 173839 284051
rect 173529 283989 173839 284023
rect 173529 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 173839 283989
rect 173529 276831 173839 283961
rect 187029 298606 187339 299134
rect 187029 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 187339 298606
rect 187029 298544 187339 298578
rect 187029 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 187339 298544
rect 187029 298482 187339 298516
rect 187029 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 187339 298482
rect 187029 298420 187339 298454
rect 187029 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 187339 298420
rect 187029 290175 187339 298392
rect 187029 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 187339 290175
rect 187029 290113 187339 290147
rect 187029 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 187339 290113
rect 187029 290051 187339 290085
rect 187029 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 187339 290051
rect 187029 289989 187339 290023
rect 187029 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 187339 289989
rect 187029 281175 187339 289961
rect 187029 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 187339 281175
rect 187029 281113 187339 281147
rect 187029 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 187339 281113
rect 187029 281051 187339 281085
rect 187029 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 187339 281051
rect 187029 280989 187339 281023
rect 187029 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 187339 280989
rect 187029 276831 187339 280961
rect 188889 299086 189199 299134
rect 188889 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 189199 299086
rect 188889 299024 189199 299058
rect 188889 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 189199 299024
rect 188889 298962 189199 298996
rect 188889 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 189199 298962
rect 188889 298900 189199 298934
rect 188889 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 189199 298900
rect 188889 293175 189199 298872
rect 188889 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 189199 293175
rect 188889 293113 189199 293147
rect 188889 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 189199 293113
rect 188889 293051 189199 293085
rect 188889 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 189199 293051
rect 188889 292989 189199 293023
rect 188889 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 189199 292989
rect 188889 284175 189199 292961
rect 188889 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 189199 284175
rect 188889 284113 189199 284147
rect 188889 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 189199 284113
rect 188889 284051 189199 284085
rect 188889 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 189199 284051
rect 188889 283989 189199 284023
rect 188889 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 189199 283989
rect 188889 276831 189199 283961
rect 202389 298606 202699 299134
rect 202389 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 202699 298606
rect 202389 298544 202699 298578
rect 202389 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 202699 298544
rect 202389 298482 202699 298516
rect 202389 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 202699 298482
rect 202389 298420 202699 298454
rect 202389 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 202699 298420
rect 202389 290175 202699 298392
rect 202389 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 202699 290175
rect 202389 290113 202699 290147
rect 202389 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 202699 290113
rect 202389 290051 202699 290085
rect 202389 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 202699 290051
rect 202389 289989 202699 290023
rect 202389 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 202699 289989
rect 202389 281175 202699 289961
rect 202389 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 202699 281175
rect 202389 281113 202699 281147
rect 202389 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 202699 281113
rect 202389 281051 202699 281085
rect 202389 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 202699 281051
rect 202389 280989 202699 281023
rect 202389 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 202699 280989
rect 202389 276831 202699 280961
rect 204249 299086 204559 299134
rect 204249 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 204559 299086
rect 204249 299024 204559 299058
rect 204249 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 204559 299024
rect 204249 298962 204559 298996
rect 204249 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 204559 298962
rect 204249 298900 204559 298934
rect 204249 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 204559 298900
rect 204249 293175 204559 298872
rect 204249 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 204559 293175
rect 204249 293113 204559 293147
rect 204249 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 204559 293113
rect 204249 293051 204559 293085
rect 204249 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 204559 293051
rect 204249 292989 204559 293023
rect 204249 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 204559 292989
rect 204249 284175 204559 292961
rect 204249 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 204559 284175
rect 204249 284113 204559 284147
rect 204249 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 204559 284113
rect 204249 284051 204559 284085
rect 204249 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 204559 284051
rect 204249 283989 204559 284023
rect 204249 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 204559 283989
rect 204249 276831 204559 283961
rect 217749 298606 218059 299134
rect 217749 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 218059 298606
rect 217749 298544 218059 298578
rect 217749 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 218059 298544
rect 217749 298482 218059 298516
rect 217749 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 218059 298482
rect 217749 298420 218059 298454
rect 217749 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 218059 298420
rect 217749 290175 218059 298392
rect 217749 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 218059 290175
rect 217749 290113 218059 290147
rect 217749 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 218059 290113
rect 217749 290051 218059 290085
rect 217749 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 218059 290051
rect 217749 289989 218059 290023
rect 217749 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 218059 289989
rect 217749 281175 218059 289961
rect 217749 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 218059 281175
rect 217749 281113 218059 281147
rect 217749 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 218059 281113
rect 217749 281051 218059 281085
rect 217749 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 218059 281051
rect 217749 280989 218059 281023
rect 217749 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 218059 280989
rect 217749 276831 218059 280961
rect 219609 299086 219919 299134
rect 219609 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 219919 299086
rect 219609 299024 219919 299058
rect 219609 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 219919 299024
rect 219609 298962 219919 298996
rect 219609 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 219919 298962
rect 219609 298900 219919 298934
rect 219609 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 219919 298900
rect 219609 293175 219919 298872
rect 219609 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 219919 293175
rect 219609 293113 219919 293147
rect 219609 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 219919 293113
rect 219609 293051 219919 293085
rect 219609 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 219919 293051
rect 219609 292989 219919 293023
rect 219609 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 219919 292989
rect 219609 284175 219919 292961
rect 219609 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 219919 284175
rect 219609 284113 219919 284147
rect 219609 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 219919 284113
rect 219609 284051 219919 284085
rect 219609 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 219919 284051
rect 219609 283989 219919 284023
rect 219609 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 219919 283989
rect 219609 276831 219919 283961
rect 233109 298606 233419 299134
rect 233109 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 233419 298606
rect 233109 298544 233419 298578
rect 233109 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 233419 298544
rect 233109 298482 233419 298516
rect 233109 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 233419 298482
rect 233109 298420 233419 298454
rect 233109 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 233419 298420
rect 233109 290175 233419 298392
rect 233109 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 233419 290175
rect 233109 290113 233419 290147
rect 233109 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 233419 290113
rect 233109 290051 233419 290085
rect 233109 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 233419 290051
rect 233109 289989 233419 290023
rect 233109 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 233419 289989
rect 233109 281175 233419 289961
rect 233109 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 233419 281175
rect 233109 281113 233419 281147
rect 233109 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 233419 281113
rect 233109 281051 233419 281085
rect 233109 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 233419 281051
rect 233109 280989 233419 281023
rect 233109 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 233419 280989
rect 233109 276831 233419 280961
rect 234969 299086 235279 299134
rect 234969 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 235279 299086
rect 234969 299024 235279 299058
rect 234969 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 235279 299024
rect 234969 298962 235279 298996
rect 234969 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 235279 298962
rect 234969 298900 235279 298934
rect 234969 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 235279 298900
rect 234969 293175 235279 298872
rect 234969 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 235279 293175
rect 234969 293113 235279 293147
rect 234969 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 235279 293113
rect 234969 293051 235279 293085
rect 234969 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 235279 293051
rect 234969 292989 235279 293023
rect 234969 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 235279 292989
rect 234969 284175 235279 292961
rect 234969 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 235279 284175
rect 234969 284113 235279 284147
rect 234969 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 235279 284113
rect 234969 284051 235279 284085
rect 234969 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 235279 284051
rect 234969 283989 235279 284023
rect 234969 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 235279 283989
rect 234969 276831 235279 283961
rect 248469 298606 248779 299134
rect 248469 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 248779 298606
rect 248469 298544 248779 298578
rect 248469 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 248779 298544
rect 248469 298482 248779 298516
rect 248469 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 248779 298482
rect 248469 298420 248779 298454
rect 248469 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 248779 298420
rect 248469 290175 248779 298392
rect 248469 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 248779 290175
rect 248469 290113 248779 290147
rect 248469 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 248779 290113
rect 248469 290051 248779 290085
rect 248469 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 248779 290051
rect 248469 289989 248779 290023
rect 248469 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 248779 289989
rect 248469 281175 248779 289961
rect 248469 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 248779 281175
rect 248469 281113 248779 281147
rect 248469 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 248779 281113
rect 248469 281051 248779 281085
rect 248469 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 248779 281051
rect 248469 280989 248779 281023
rect 248469 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 248779 280989
rect 248469 276831 248779 280961
rect 250329 299086 250639 299134
rect 250329 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 250639 299086
rect 250329 299024 250639 299058
rect 250329 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 250639 299024
rect 250329 298962 250639 298996
rect 250329 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 250639 298962
rect 250329 298900 250639 298934
rect 250329 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 250639 298900
rect 250329 293175 250639 298872
rect 250329 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 250639 293175
rect 250329 293113 250639 293147
rect 250329 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 250639 293113
rect 250329 293051 250639 293085
rect 250329 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 250639 293051
rect 250329 292989 250639 293023
rect 250329 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 250639 292989
rect 250329 284175 250639 292961
rect 250329 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 250639 284175
rect 250329 284113 250639 284147
rect 250329 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 250639 284113
rect 250329 284051 250639 284085
rect 250329 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 250639 284051
rect 250329 283989 250639 284023
rect 250329 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 250639 283989
rect 250329 276831 250639 283961
rect 263829 298606 264139 299134
rect 263829 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 264139 298606
rect 263829 298544 264139 298578
rect 263829 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 264139 298544
rect 263829 298482 264139 298516
rect 263829 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 264139 298482
rect 263829 298420 264139 298454
rect 263829 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 264139 298420
rect 263829 290175 264139 298392
rect 263829 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 264139 290175
rect 263829 290113 264139 290147
rect 263829 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 264139 290113
rect 263829 290051 264139 290085
rect 263829 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 264139 290051
rect 263829 289989 264139 290023
rect 263829 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 264139 289989
rect 263829 281175 264139 289961
rect 263829 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 264139 281175
rect 263829 281113 264139 281147
rect 263829 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 264139 281113
rect 263829 281051 264139 281085
rect 263829 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 264139 281051
rect 263829 280989 264139 281023
rect 263829 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 264139 280989
rect 263829 276831 264139 280961
rect 265689 299086 265999 299134
rect 265689 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 265999 299086
rect 265689 299024 265999 299058
rect 265689 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 265999 299024
rect 265689 298962 265999 298996
rect 265689 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 265999 298962
rect 265689 298900 265999 298934
rect 265689 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 265999 298900
rect 265689 293175 265999 298872
rect 265689 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 265999 293175
rect 265689 293113 265999 293147
rect 265689 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 265999 293113
rect 265689 293051 265999 293085
rect 265689 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 265999 293051
rect 265689 292989 265999 293023
rect 265689 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 265999 292989
rect 265689 284175 265999 292961
rect 265689 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 265999 284175
rect 265689 284113 265999 284147
rect 265689 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 265999 284113
rect 265689 284051 265999 284085
rect 265689 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 265999 284051
rect 265689 283989 265999 284023
rect 265689 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 265999 283989
rect 265689 276831 265999 283961
rect 279189 298606 279499 299134
rect 279189 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 279499 298606
rect 279189 298544 279499 298578
rect 279189 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 279499 298544
rect 279189 298482 279499 298516
rect 279189 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 279499 298482
rect 279189 298420 279499 298454
rect 279189 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 279499 298420
rect 279189 290175 279499 298392
rect 279189 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 279499 290175
rect 279189 290113 279499 290147
rect 279189 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 279499 290113
rect 279189 290051 279499 290085
rect 279189 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 279499 290051
rect 279189 289989 279499 290023
rect 279189 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 279499 289989
rect 279189 281175 279499 289961
rect 279189 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 279499 281175
rect 279189 281113 279499 281147
rect 279189 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 279499 281113
rect 279189 281051 279499 281085
rect 279189 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 279499 281051
rect 279189 280989 279499 281023
rect 279189 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 279499 280989
rect 96729 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 97039 275175
rect 96729 275113 97039 275147
rect 96729 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 97039 275113
rect 96729 275051 97039 275085
rect 96729 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 97039 275051
rect 96729 274989 97039 275023
rect 109904 275175 110064 275192
rect 109904 275147 109939 275175
rect 109967 275147 110001 275175
rect 110029 275147 110064 275175
rect 109904 275113 110064 275147
rect 109904 275085 109939 275113
rect 109967 275085 110001 275113
rect 110029 275085 110064 275113
rect 109904 275051 110064 275085
rect 109904 275023 109939 275051
rect 109967 275023 110001 275051
rect 110029 275023 110064 275051
rect 96729 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 97039 274989
rect 96729 266175 97039 274961
rect 96729 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 97039 266175
rect 96729 266113 97039 266147
rect 96729 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 97039 266113
rect 96729 266051 97039 266085
rect 96729 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 97039 266051
rect 96729 265989 97039 266023
rect 96729 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 97039 265989
rect 96729 257175 97039 265961
rect 96729 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 97039 257175
rect 96729 257113 97039 257147
rect 96729 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 97039 257113
rect 96729 257051 97039 257085
rect 96729 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 97039 257051
rect 96729 256989 97039 257023
rect 96729 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 97039 256989
rect 96729 248175 97039 256961
rect 96729 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 97039 248175
rect 96729 248113 97039 248147
rect 96729 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 97039 248113
rect 96729 248051 97039 248085
rect 96729 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 97039 248051
rect 96729 247989 97039 248023
rect 96729 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 97039 247989
rect 96729 239175 97039 247961
rect 96729 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 97039 239175
rect 96729 239113 97039 239147
rect 96729 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 97039 239113
rect 96729 239051 97039 239085
rect 96729 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 97039 239051
rect 96729 238989 97039 239023
rect 96729 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 97039 238989
rect 96729 230175 97039 238961
rect 96729 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 97039 230175
rect 96729 230113 97039 230147
rect 96729 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 97039 230113
rect 96729 230051 97039 230085
rect 96729 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 97039 230051
rect 96729 229989 97039 230023
rect 96729 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 97039 229989
rect 96729 221175 97039 229961
rect 96729 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 97039 221175
rect 96729 221113 97039 221147
rect 96729 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 97039 221113
rect 96729 221051 97039 221085
rect 96729 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 97039 221051
rect 96729 220989 97039 221023
rect 96729 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 97039 220989
rect 96729 212175 97039 220961
rect 96729 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 97039 212175
rect 96729 212113 97039 212147
rect 96729 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 97039 212113
rect 96729 212051 97039 212085
rect 96729 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 97039 212051
rect 96729 211989 97039 212023
rect 96729 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 97039 211989
rect 96729 203175 97039 211961
rect 96729 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 97039 203175
rect 96729 203113 97039 203147
rect 96729 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 97039 203113
rect 96729 203051 97039 203085
rect 96729 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 97039 203051
rect 96729 202989 97039 203023
rect 96729 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 97039 202989
rect 96729 194175 97039 202961
rect 96729 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 97039 194175
rect 96729 194113 97039 194147
rect 96729 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 97039 194113
rect 96729 194051 97039 194085
rect 96729 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 97039 194051
rect 96729 193989 97039 194023
rect 96729 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 97039 193989
rect 96729 185175 97039 193961
rect 98686 275002 98714 275007
rect 96729 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 97039 185175
rect 96729 185113 97039 185147
rect 96729 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 97039 185113
rect 96729 185051 97039 185085
rect 96729 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 97039 185051
rect 96729 184989 97039 185023
rect 96729 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 97039 184989
rect 96729 176175 97039 184961
rect 96729 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 97039 176175
rect 96729 176113 97039 176147
rect 96729 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 97039 176113
rect 96729 176051 97039 176085
rect 96729 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 97039 176051
rect 96729 175989 97039 176023
rect 96729 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 97039 175989
rect 96729 167175 97039 175961
rect 96729 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 97039 167175
rect 96729 167113 97039 167147
rect 96729 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 97039 167113
rect 96729 167051 97039 167085
rect 96729 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 97039 167051
rect 96729 166989 97039 167023
rect 96729 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 97039 166989
rect 96729 158175 97039 166961
rect 96729 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 97039 158175
rect 96729 158113 97039 158147
rect 96729 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 97039 158113
rect 96729 158051 97039 158085
rect 96729 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 97039 158051
rect 96729 157989 97039 158023
rect 96729 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 97039 157989
rect 96729 149175 97039 157961
rect 96729 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 97039 149175
rect 96729 149113 97039 149147
rect 96729 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 97039 149113
rect 96729 149051 97039 149085
rect 96729 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 97039 149051
rect 96729 148989 97039 149023
rect 96729 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 97039 148989
rect 96729 140175 97039 148961
rect 96729 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 97039 140175
rect 96729 140113 97039 140147
rect 96729 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 97039 140113
rect 96729 140051 97039 140085
rect 96729 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 97039 140051
rect 96729 139989 97039 140023
rect 96729 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 97039 139989
rect 96729 131175 97039 139961
rect 96729 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 97039 131175
rect 96729 131113 97039 131147
rect 96729 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 97039 131113
rect 96729 131051 97039 131085
rect 96729 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 97039 131051
rect 96729 130989 97039 131023
rect 96729 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130961 97039 130989
rect 96729 122175 97039 130961
rect 96729 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 97039 122175
rect 96729 122113 97039 122147
rect 96729 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 97039 122113
rect 96729 122051 97039 122085
rect 96729 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 97039 122051
rect 96729 121989 97039 122023
rect 96729 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 97039 121989
rect 96729 113175 97039 121961
rect 96729 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 97039 113175
rect 96729 113113 97039 113147
rect 96729 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 97039 113113
rect 96729 113051 97039 113085
rect 96729 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 97039 113051
rect 96729 112989 97039 113023
rect 96729 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 97039 112989
rect 96729 104175 97039 112961
rect 96729 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 97039 104175
rect 96729 104113 97039 104147
rect 96729 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 97039 104113
rect 96729 104051 97039 104085
rect 96729 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 97039 104051
rect 96729 103989 97039 104023
rect 96729 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 97039 103989
rect 96729 95175 97039 103961
rect 96729 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 97039 95175
rect 96729 95113 97039 95147
rect 96729 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 97039 95113
rect 96729 95051 97039 95085
rect 96729 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 97039 95051
rect 96729 94989 97039 95023
rect 96729 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 97039 94989
rect 96729 86175 97039 94961
rect 96729 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 97039 86175
rect 96729 86113 97039 86147
rect 96729 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 97039 86113
rect 96729 86051 97039 86085
rect 96729 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 97039 86051
rect 96729 85989 97039 86023
rect 96729 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 97039 85989
rect 96729 77175 97039 85961
rect 98630 186298 98658 186303
rect 98630 81914 98658 186270
rect 98686 166586 98714 274974
rect 109904 274989 110064 275023
rect 109904 274961 109939 274989
rect 109967 274961 110001 274989
rect 110029 274961 110064 274989
rect 109904 274944 110064 274961
rect 125264 275175 125424 275192
rect 125264 275147 125299 275175
rect 125327 275147 125361 275175
rect 125389 275147 125424 275175
rect 125264 275113 125424 275147
rect 125264 275085 125299 275113
rect 125327 275085 125361 275113
rect 125389 275085 125424 275113
rect 125264 275051 125424 275085
rect 125264 275023 125299 275051
rect 125327 275023 125361 275051
rect 125389 275023 125424 275051
rect 125264 274989 125424 275023
rect 125264 274961 125299 274989
rect 125327 274961 125361 274989
rect 125389 274961 125424 274989
rect 125264 274944 125424 274961
rect 140624 275175 140784 275192
rect 140624 275147 140659 275175
rect 140687 275147 140721 275175
rect 140749 275147 140784 275175
rect 140624 275113 140784 275147
rect 140624 275085 140659 275113
rect 140687 275085 140721 275113
rect 140749 275085 140784 275113
rect 140624 275051 140784 275085
rect 140624 275023 140659 275051
rect 140687 275023 140721 275051
rect 140749 275023 140784 275051
rect 140624 274989 140784 275023
rect 140624 274961 140659 274989
rect 140687 274961 140721 274989
rect 140749 274961 140784 274989
rect 140624 274944 140784 274961
rect 155984 275175 156144 275192
rect 155984 275147 156019 275175
rect 156047 275147 156081 275175
rect 156109 275147 156144 275175
rect 155984 275113 156144 275147
rect 155984 275085 156019 275113
rect 156047 275085 156081 275113
rect 156109 275085 156144 275113
rect 155984 275051 156144 275085
rect 155984 275023 156019 275051
rect 156047 275023 156081 275051
rect 156109 275023 156144 275051
rect 155984 274989 156144 275023
rect 155984 274961 156019 274989
rect 156047 274961 156081 274989
rect 156109 274961 156144 274989
rect 155984 274944 156144 274961
rect 171344 275175 171504 275192
rect 171344 275147 171379 275175
rect 171407 275147 171441 275175
rect 171469 275147 171504 275175
rect 171344 275113 171504 275147
rect 171344 275085 171379 275113
rect 171407 275085 171441 275113
rect 171469 275085 171504 275113
rect 171344 275051 171504 275085
rect 171344 275023 171379 275051
rect 171407 275023 171441 275051
rect 171469 275023 171504 275051
rect 171344 274989 171504 275023
rect 171344 274961 171379 274989
rect 171407 274961 171441 274989
rect 171469 274961 171504 274989
rect 171344 274944 171504 274961
rect 186704 275175 186864 275192
rect 186704 275147 186739 275175
rect 186767 275147 186801 275175
rect 186829 275147 186864 275175
rect 186704 275113 186864 275147
rect 186704 275085 186739 275113
rect 186767 275085 186801 275113
rect 186829 275085 186864 275113
rect 186704 275051 186864 275085
rect 186704 275023 186739 275051
rect 186767 275023 186801 275051
rect 186829 275023 186864 275051
rect 186704 274989 186864 275023
rect 186704 274961 186739 274989
rect 186767 274961 186801 274989
rect 186829 274961 186864 274989
rect 186704 274944 186864 274961
rect 202064 275175 202224 275192
rect 202064 275147 202099 275175
rect 202127 275147 202161 275175
rect 202189 275147 202224 275175
rect 202064 275113 202224 275147
rect 202064 275085 202099 275113
rect 202127 275085 202161 275113
rect 202189 275085 202224 275113
rect 202064 275051 202224 275085
rect 202064 275023 202099 275051
rect 202127 275023 202161 275051
rect 202189 275023 202224 275051
rect 202064 274989 202224 275023
rect 202064 274961 202099 274989
rect 202127 274961 202161 274989
rect 202189 274961 202224 274989
rect 202064 274944 202224 274961
rect 217424 275175 217584 275192
rect 217424 275147 217459 275175
rect 217487 275147 217521 275175
rect 217549 275147 217584 275175
rect 217424 275113 217584 275147
rect 217424 275085 217459 275113
rect 217487 275085 217521 275113
rect 217549 275085 217584 275113
rect 217424 275051 217584 275085
rect 217424 275023 217459 275051
rect 217487 275023 217521 275051
rect 217549 275023 217584 275051
rect 217424 274989 217584 275023
rect 217424 274961 217459 274989
rect 217487 274961 217521 274989
rect 217549 274961 217584 274989
rect 217424 274944 217584 274961
rect 232784 275175 232944 275192
rect 232784 275147 232819 275175
rect 232847 275147 232881 275175
rect 232909 275147 232944 275175
rect 232784 275113 232944 275147
rect 232784 275085 232819 275113
rect 232847 275085 232881 275113
rect 232909 275085 232944 275113
rect 232784 275051 232944 275085
rect 232784 275023 232819 275051
rect 232847 275023 232881 275051
rect 232909 275023 232944 275051
rect 232784 274989 232944 275023
rect 232784 274961 232819 274989
rect 232847 274961 232881 274989
rect 232909 274961 232944 274989
rect 232784 274944 232944 274961
rect 248144 275175 248304 275192
rect 248144 275147 248179 275175
rect 248207 275147 248241 275175
rect 248269 275147 248304 275175
rect 248144 275113 248304 275147
rect 248144 275085 248179 275113
rect 248207 275085 248241 275113
rect 248269 275085 248304 275113
rect 248144 275051 248304 275085
rect 248144 275023 248179 275051
rect 248207 275023 248241 275051
rect 248269 275023 248304 275051
rect 248144 274989 248304 275023
rect 248144 274961 248179 274989
rect 248207 274961 248241 274989
rect 248269 274961 248304 274989
rect 248144 274944 248304 274961
rect 263504 275175 263664 275192
rect 263504 275147 263539 275175
rect 263567 275147 263601 275175
rect 263629 275147 263664 275175
rect 263504 275113 263664 275147
rect 263504 275085 263539 275113
rect 263567 275085 263601 275113
rect 263629 275085 263664 275113
rect 263504 275051 263664 275085
rect 263504 275023 263539 275051
rect 263567 275023 263601 275051
rect 263629 275023 263664 275051
rect 263504 274989 263664 275023
rect 263504 274961 263539 274989
rect 263567 274961 263601 274989
rect 263629 274961 263664 274989
rect 263504 274944 263664 274961
rect 278864 275175 279024 275192
rect 278864 275147 278899 275175
rect 278927 275147 278961 275175
rect 278989 275147 279024 275175
rect 278864 275113 279024 275147
rect 278864 275085 278899 275113
rect 278927 275085 278961 275113
rect 278989 275085 279024 275113
rect 278864 275051 279024 275085
rect 278864 275023 278899 275051
rect 278927 275023 278961 275051
rect 278989 275023 279024 275051
rect 278864 274989 279024 275023
rect 278864 274961 278899 274989
rect 278927 274961 278961 274989
rect 278989 274961 279024 274989
rect 278864 274944 279024 274961
rect 102224 272175 102384 272192
rect 102224 272147 102259 272175
rect 102287 272147 102321 272175
rect 102349 272147 102384 272175
rect 102224 272113 102384 272147
rect 102224 272085 102259 272113
rect 102287 272085 102321 272113
rect 102349 272085 102384 272113
rect 102224 272051 102384 272085
rect 102224 272023 102259 272051
rect 102287 272023 102321 272051
rect 102349 272023 102384 272051
rect 102224 271989 102384 272023
rect 102224 271961 102259 271989
rect 102287 271961 102321 271989
rect 102349 271961 102384 271989
rect 102224 271944 102384 271961
rect 117584 272175 117744 272192
rect 117584 272147 117619 272175
rect 117647 272147 117681 272175
rect 117709 272147 117744 272175
rect 117584 272113 117744 272147
rect 117584 272085 117619 272113
rect 117647 272085 117681 272113
rect 117709 272085 117744 272113
rect 117584 272051 117744 272085
rect 117584 272023 117619 272051
rect 117647 272023 117681 272051
rect 117709 272023 117744 272051
rect 117584 271989 117744 272023
rect 117584 271961 117619 271989
rect 117647 271961 117681 271989
rect 117709 271961 117744 271989
rect 117584 271944 117744 271961
rect 132944 272175 133104 272192
rect 132944 272147 132979 272175
rect 133007 272147 133041 272175
rect 133069 272147 133104 272175
rect 132944 272113 133104 272147
rect 132944 272085 132979 272113
rect 133007 272085 133041 272113
rect 133069 272085 133104 272113
rect 132944 272051 133104 272085
rect 132944 272023 132979 272051
rect 133007 272023 133041 272051
rect 133069 272023 133104 272051
rect 132944 271989 133104 272023
rect 132944 271961 132979 271989
rect 133007 271961 133041 271989
rect 133069 271961 133104 271989
rect 132944 271944 133104 271961
rect 148304 272175 148464 272192
rect 148304 272147 148339 272175
rect 148367 272147 148401 272175
rect 148429 272147 148464 272175
rect 148304 272113 148464 272147
rect 148304 272085 148339 272113
rect 148367 272085 148401 272113
rect 148429 272085 148464 272113
rect 148304 272051 148464 272085
rect 148304 272023 148339 272051
rect 148367 272023 148401 272051
rect 148429 272023 148464 272051
rect 148304 271989 148464 272023
rect 148304 271961 148339 271989
rect 148367 271961 148401 271989
rect 148429 271961 148464 271989
rect 148304 271944 148464 271961
rect 163664 272175 163824 272192
rect 163664 272147 163699 272175
rect 163727 272147 163761 272175
rect 163789 272147 163824 272175
rect 163664 272113 163824 272147
rect 163664 272085 163699 272113
rect 163727 272085 163761 272113
rect 163789 272085 163824 272113
rect 163664 272051 163824 272085
rect 163664 272023 163699 272051
rect 163727 272023 163761 272051
rect 163789 272023 163824 272051
rect 163664 271989 163824 272023
rect 163664 271961 163699 271989
rect 163727 271961 163761 271989
rect 163789 271961 163824 271989
rect 163664 271944 163824 271961
rect 179024 272175 179184 272192
rect 179024 272147 179059 272175
rect 179087 272147 179121 272175
rect 179149 272147 179184 272175
rect 179024 272113 179184 272147
rect 179024 272085 179059 272113
rect 179087 272085 179121 272113
rect 179149 272085 179184 272113
rect 179024 272051 179184 272085
rect 179024 272023 179059 272051
rect 179087 272023 179121 272051
rect 179149 272023 179184 272051
rect 179024 271989 179184 272023
rect 179024 271961 179059 271989
rect 179087 271961 179121 271989
rect 179149 271961 179184 271989
rect 179024 271944 179184 271961
rect 194384 272175 194544 272192
rect 194384 272147 194419 272175
rect 194447 272147 194481 272175
rect 194509 272147 194544 272175
rect 194384 272113 194544 272147
rect 194384 272085 194419 272113
rect 194447 272085 194481 272113
rect 194509 272085 194544 272113
rect 194384 272051 194544 272085
rect 194384 272023 194419 272051
rect 194447 272023 194481 272051
rect 194509 272023 194544 272051
rect 194384 271989 194544 272023
rect 194384 271961 194419 271989
rect 194447 271961 194481 271989
rect 194509 271961 194544 271989
rect 194384 271944 194544 271961
rect 209744 272175 209904 272192
rect 209744 272147 209779 272175
rect 209807 272147 209841 272175
rect 209869 272147 209904 272175
rect 209744 272113 209904 272147
rect 209744 272085 209779 272113
rect 209807 272085 209841 272113
rect 209869 272085 209904 272113
rect 209744 272051 209904 272085
rect 209744 272023 209779 272051
rect 209807 272023 209841 272051
rect 209869 272023 209904 272051
rect 209744 271989 209904 272023
rect 209744 271961 209779 271989
rect 209807 271961 209841 271989
rect 209869 271961 209904 271989
rect 209744 271944 209904 271961
rect 225104 272175 225264 272192
rect 225104 272147 225139 272175
rect 225167 272147 225201 272175
rect 225229 272147 225264 272175
rect 225104 272113 225264 272147
rect 225104 272085 225139 272113
rect 225167 272085 225201 272113
rect 225229 272085 225264 272113
rect 225104 272051 225264 272085
rect 225104 272023 225139 272051
rect 225167 272023 225201 272051
rect 225229 272023 225264 272051
rect 225104 271989 225264 272023
rect 225104 271961 225139 271989
rect 225167 271961 225201 271989
rect 225229 271961 225264 271989
rect 225104 271944 225264 271961
rect 240464 272175 240624 272192
rect 240464 272147 240499 272175
rect 240527 272147 240561 272175
rect 240589 272147 240624 272175
rect 240464 272113 240624 272147
rect 240464 272085 240499 272113
rect 240527 272085 240561 272113
rect 240589 272085 240624 272113
rect 240464 272051 240624 272085
rect 240464 272023 240499 272051
rect 240527 272023 240561 272051
rect 240589 272023 240624 272051
rect 240464 271989 240624 272023
rect 240464 271961 240499 271989
rect 240527 271961 240561 271989
rect 240589 271961 240624 271989
rect 240464 271944 240624 271961
rect 255824 272175 255984 272192
rect 255824 272147 255859 272175
rect 255887 272147 255921 272175
rect 255949 272147 255984 272175
rect 255824 272113 255984 272147
rect 255824 272085 255859 272113
rect 255887 272085 255921 272113
rect 255949 272085 255984 272113
rect 255824 272051 255984 272085
rect 255824 272023 255859 272051
rect 255887 272023 255921 272051
rect 255949 272023 255984 272051
rect 255824 271989 255984 272023
rect 255824 271961 255859 271989
rect 255887 271961 255921 271989
rect 255949 271961 255984 271989
rect 255824 271944 255984 271961
rect 271184 272175 271344 272192
rect 271184 272147 271219 272175
rect 271247 272147 271281 272175
rect 271309 272147 271344 272175
rect 271184 272113 271344 272147
rect 271184 272085 271219 272113
rect 271247 272085 271281 272113
rect 271309 272085 271344 272113
rect 271184 272051 271344 272085
rect 271184 272023 271219 272051
rect 271247 272023 271281 272051
rect 271309 272023 271344 272051
rect 271184 271989 271344 272023
rect 271184 271961 271219 271989
rect 271247 271961 271281 271989
rect 271309 271961 271344 271989
rect 271184 271944 271344 271961
rect 279189 272175 279499 280961
rect 279189 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 279499 272175
rect 279189 272113 279499 272147
rect 279189 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 279499 272113
rect 279189 272051 279499 272085
rect 279189 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 279499 272051
rect 279189 271989 279499 272023
rect 279189 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 279499 271989
rect 109904 266175 110064 266192
rect 109904 266147 109939 266175
rect 109967 266147 110001 266175
rect 110029 266147 110064 266175
rect 109904 266113 110064 266147
rect 109904 266085 109939 266113
rect 109967 266085 110001 266113
rect 110029 266085 110064 266113
rect 109904 266051 110064 266085
rect 109904 266023 109939 266051
rect 109967 266023 110001 266051
rect 110029 266023 110064 266051
rect 109904 265989 110064 266023
rect 109904 265961 109939 265989
rect 109967 265961 110001 265989
rect 110029 265961 110064 265989
rect 109904 265944 110064 265961
rect 125264 266175 125424 266192
rect 125264 266147 125299 266175
rect 125327 266147 125361 266175
rect 125389 266147 125424 266175
rect 125264 266113 125424 266147
rect 125264 266085 125299 266113
rect 125327 266085 125361 266113
rect 125389 266085 125424 266113
rect 125264 266051 125424 266085
rect 125264 266023 125299 266051
rect 125327 266023 125361 266051
rect 125389 266023 125424 266051
rect 125264 265989 125424 266023
rect 125264 265961 125299 265989
rect 125327 265961 125361 265989
rect 125389 265961 125424 265989
rect 125264 265944 125424 265961
rect 140624 266175 140784 266192
rect 140624 266147 140659 266175
rect 140687 266147 140721 266175
rect 140749 266147 140784 266175
rect 140624 266113 140784 266147
rect 140624 266085 140659 266113
rect 140687 266085 140721 266113
rect 140749 266085 140784 266113
rect 140624 266051 140784 266085
rect 140624 266023 140659 266051
rect 140687 266023 140721 266051
rect 140749 266023 140784 266051
rect 140624 265989 140784 266023
rect 140624 265961 140659 265989
rect 140687 265961 140721 265989
rect 140749 265961 140784 265989
rect 140624 265944 140784 265961
rect 155984 266175 156144 266192
rect 155984 266147 156019 266175
rect 156047 266147 156081 266175
rect 156109 266147 156144 266175
rect 155984 266113 156144 266147
rect 155984 266085 156019 266113
rect 156047 266085 156081 266113
rect 156109 266085 156144 266113
rect 155984 266051 156144 266085
rect 155984 266023 156019 266051
rect 156047 266023 156081 266051
rect 156109 266023 156144 266051
rect 155984 265989 156144 266023
rect 155984 265961 156019 265989
rect 156047 265961 156081 265989
rect 156109 265961 156144 265989
rect 155984 265944 156144 265961
rect 171344 266175 171504 266192
rect 171344 266147 171379 266175
rect 171407 266147 171441 266175
rect 171469 266147 171504 266175
rect 171344 266113 171504 266147
rect 171344 266085 171379 266113
rect 171407 266085 171441 266113
rect 171469 266085 171504 266113
rect 171344 266051 171504 266085
rect 171344 266023 171379 266051
rect 171407 266023 171441 266051
rect 171469 266023 171504 266051
rect 171344 265989 171504 266023
rect 171344 265961 171379 265989
rect 171407 265961 171441 265989
rect 171469 265961 171504 265989
rect 171344 265944 171504 265961
rect 186704 266175 186864 266192
rect 186704 266147 186739 266175
rect 186767 266147 186801 266175
rect 186829 266147 186864 266175
rect 186704 266113 186864 266147
rect 186704 266085 186739 266113
rect 186767 266085 186801 266113
rect 186829 266085 186864 266113
rect 186704 266051 186864 266085
rect 186704 266023 186739 266051
rect 186767 266023 186801 266051
rect 186829 266023 186864 266051
rect 186704 265989 186864 266023
rect 186704 265961 186739 265989
rect 186767 265961 186801 265989
rect 186829 265961 186864 265989
rect 186704 265944 186864 265961
rect 202064 266175 202224 266192
rect 202064 266147 202099 266175
rect 202127 266147 202161 266175
rect 202189 266147 202224 266175
rect 202064 266113 202224 266147
rect 202064 266085 202099 266113
rect 202127 266085 202161 266113
rect 202189 266085 202224 266113
rect 202064 266051 202224 266085
rect 202064 266023 202099 266051
rect 202127 266023 202161 266051
rect 202189 266023 202224 266051
rect 202064 265989 202224 266023
rect 202064 265961 202099 265989
rect 202127 265961 202161 265989
rect 202189 265961 202224 265989
rect 202064 265944 202224 265961
rect 217424 266175 217584 266192
rect 217424 266147 217459 266175
rect 217487 266147 217521 266175
rect 217549 266147 217584 266175
rect 217424 266113 217584 266147
rect 217424 266085 217459 266113
rect 217487 266085 217521 266113
rect 217549 266085 217584 266113
rect 217424 266051 217584 266085
rect 217424 266023 217459 266051
rect 217487 266023 217521 266051
rect 217549 266023 217584 266051
rect 217424 265989 217584 266023
rect 217424 265961 217459 265989
rect 217487 265961 217521 265989
rect 217549 265961 217584 265989
rect 217424 265944 217584 265961
rect 232784 266175 232944 266192
rect 232784 266147 232819 266175
rect 232847 266147 232881 266175
rect 232909 266147 232944 266175
rect 232784 266113 232944 266147
rect 232784 266085 232819 266113
rect 232847 266085 232881 266113
rect 232909 266085 232944 266113
rect 232784 266051 232944 266085
rect 232784 266023 232819 266051
rect 232847 266023 232881 266051
rect 232909 266023 232944 266051
rect 232784 265989 232944 266023
rect 232784 265961 232819 265989
rect 232847 265961 232881 265989
rect 232909 265961 232944 265989
rect 232784 265944 232944 265961
rect 248144 266175 248304 266192
rect 248144 266147 248179 266175
rect 248207 266147 248241 266175
rect 248269 266147 248304 266175
rect 248144 266113 248304 266147
rect 248144 266085 248179 266113
rect 248207 266085 248241 266113
rect 248269 266085 248304 266113
rect 248144 266051 248304 266085
rect 248144 266023 248179 266051
rect 248207 266023 248241 266051
rect 248269 266023 248304 266051
rect 248144 265989 248304 266023
rect 248144 265961 248179 265989
rect 248207 265961 248241 265989
rect 248269 265961 248304 265989
rect 248144 265944 248304 265961
rect 263504 266175 263664 266192
rect 263504 266147 263539 266175
rect 263567 266147 263601 266175
rect 263629 266147 263664 266175
rect 263504 266113 263664 266147
rect 263504 266085 263539 266113
rect 263567 266085 263601 266113
rect 263629 266085 263664 266113
rect 263504 266051 263664 266085
rect 263504 266023 263539 266051
rect 263567 266023 263601 266051
rect 263629 266023 263664 266051
rect 263504 265989 263664 266023
rect 263504 265961 263539 265989
rect 263567 265961 263601 265989
rect 263629 265961 263664 265989
rect 263504 265944 263664 265961
rect 278864 266175 279024 266192
rect 278864 266147 278899 266175
rect 278927 266147 278961 266175
rect 278989 266147 279024 266175
rect 278864 266113 279024 266147
rect 278864 266085 278899 266113
rect 278927 266085 278961 266113
rect 278989 266085 279024 266113
rect 278864 266051 279024 266085
rect 278864 266023 278899 266051
rect 278927 266023 278961 266051
rect 278989 266023 279024 266051
rect 278864 265989 279024 266023
rect 278864 265961 278899 265989
rect 278927 265961 278961 265989
rect 278989 265961 279024 265989
rect 278864 265944 279024 265961
rect 102224 263175 102384 263192
rect 102224 263147 102259 263175
rect 102287 263147 102321 263175
rect 102349 263147 102384 263175
rect 102224 263113 102384 263147
rect 102224 263085 102259 263113
rect 102287 263085 102321 263113
rect 102349 263085 102384 263113
rect 102224 263051 102384 263085
rect 102224 263023 102259 263051
rect 102287 263023 102321 263051
rect 102349 263023 102384 263051
rect 102224 262989 102384 263023
rect 102224 262961 102259 262989
rect 102287 262961 102321 262989
rect 102349 262961 102384 262989
rect 102224 262944 102384 262961
rect 117584 263175 117744 263192
rect 117584 263147 117619 263175
rect 117647 263147 117681 263175
rect 117709 263147 117744 263175
rect 117584 263113 117744 263147
rect 117584 263085 117619 263113
rect 117647 263085 117681 263113
rect 117709 263085 117744 263113
rect 117584 263051 117744 263085
rect 117584 263023 117619 263051
rect 117647 263023 117681 263051
rect 117709 263023 117744 263051
rect 117584 262989 117744 263023
rect 117584 262961 117619 262989
rect 117647 262961 117681 262989
rect 117709 262961 117744 262989
rect 117584 262944 117744 262961
rect 132944 263175 133104 263192
rect 132944 263147 132979 263175
rect 133007 263147 133041 263175
rect 133069 263147 133104 263175
rect 132944 263113 133104 263147
rect 132944 263085 132979 263113
rect 133007 263085 133041 263113
rect 133069 263085 133104 263113
rect 132944 263051 133104 263085
rect 132944 263023 132979 263051
rect 133007 263023 133041 263051
rect 133069 263023 133104 263051
rect 132944 262989 133104 263023
rect 132944 262961 132979 262989
rect 133007 262961 133041 262989
rect 133069 262961 133104 262989
rect 132944 262944 133104 262961
rect 148304 263175 148464 263192
rect 148304 263147 148339 263175
rect 148367 263147 148401 263175
rect 148429 263147 148464 263175
rect 148304 263113 148464 263147
rect 148304 263085 148339 263113
rect 148367 263085 148401 263113
rect 148429 263085 148464 263113
rect 148304 263051 148464 263085
rect 148304 263023 148339 263051
rect 148367 263023 148401 263051
rect 148429 263023 148464 263051
rect 148304 262989 148464 263023
rect 148304 262961 148339 262989
rect 148367 262961 148401 262989
rect 148429 262961 148464 262989
rect 148304 262944 148464 262961
rect 163664 263175 163824 263192
rect 163664 263147 163699 263175
rect 163727 263147 163761 263175
rect 163789 263147 163824 263175
rect 163664 263113 163824 263147
rect 163664 263085 163699 263113
rect 163727 263085 163761 263113
rect 163789 263085 163824 263113
rect 163664 263051 163824 263085
rect 163664 263023 163699 263051
rect 163727 263023 163761 263051
rect 163789 263023 163824 263051
rect 163664 262989 163824 263023
rect 163664 262961 163699 262989
rect 163727 262961 163761 262989
rect 163789 262961 163824 262989
rect 163664 262944 163824 262961
rect 179024 263175 179184 263192
rect 179024 263147 179059 263175
rect 179087 263147 179121 263175
rect 179149 263147 179184 263175
rect 179024 263113 179184 263147
rect 179024 263085 179059 263113
rect 179087 263085 179121 263113
rect 179149 263085 179184 263113
rect 179024 263051 179184 263085
rect 179024 263023 179059 263051
rect 179087 263023 179121 263051
rect 179149 263023 179184 263051
rect 179024 262989 179184 263023
rect 179024 262961 179059 262989
rect 179087 262961 179121 262989
rect 179149 262961 179184 262989
rect 179024 262944 179184 262961
rect 194384 263175 194544 263192
rect 194384 263147 194419 263175
rect 194447 263147 194481 263175
rect 194509 263147 194544 263175
rect 194384 263113 194544 263147
rect 194384 263085 194419 263113
rect 194447 263085 194481 263113
rect 194509 263085 194544 263113
rect 194384 263051 194544 263085
rect 194384 263023 194419 263051
rect 194447 263023 194481 263051
rect 194509 263023 194544 263051
rect 194384 262989 194544 263023
rect 194384 262961 194419 262989
rect 194447 262961 194481 262989
rect 194509 262961 194544 262989
rect 194384 262944 194544 262961
rect 209744 263175 209904 263192
rect 209744 263147 209779 263175
rect 209807 263147 209841 263175
rect 209869 263147 209904 263175
rect 209744 263113 209904 263147
rect 209744 263085 209779 263113
rect 209807 263085 209841 263113
rect 209869 263085 209904 263113
rect 209744 263051 209904 263085
rect 209744 263023 209779 263051
rect 209807 263023 209841 263051
rect 209869 263023 209904 263051
rect 209744 262989 209904 263023
rect 209744 262961 209779 262989
rect 209807 262961 209841 262989
rect 209869 262961 209904 262989
rect 209744 262944 209904 262961
rect 225104 263175 225264 263192
rect 225104 263147 225139 263175
rect 225167 263147 225201 263175
rect 225229 263147 225264 263175
rect 225104 263113 225264 263147
rect 225104 263085 225139 263113
rect 225167 263085 225201 263113
rect 225229 263085 225264 263113
rect 225104 263051 225264 263085
rect 225104 263023 225139 263051
rect 225167 263023 225201 263051
rect 225229 263023 225264 263051
rect 225104 262989 225264 263023
rect 225104 262961 225139 262989
rect 225167 262961 225201 262989
rect 225229 262961 225264 262989
rect 225104 262944 225264 262961
rect 240464 263175 240624 263192
rect 240464 263147 240499 263175
rect 240527 263147 240561 263175
rect 240589 263147 240624 263175
rect 240464 263113 240624 263147
rect 240464 263085 240499 263113
rect 240527 263085 240561 263113
rect 240589 263085 240624 263113
rect 240464 263051 240624 263085
rect 240464 263023 240499 263051
rect 240527 263023 240561 263051
rect 240589 263023 240624 263051
rect 240464 262989 240624 263023
rect 240464 262961 240499 262989
rect 240527 262961 240561 262989
rect 240589 262961 240624 262989
rect 240464 262944 240624 262961
rect 255824 263175 255984 263192
rect 255824 263147 255859 263175
rect 255887 263147 255921 263175
rect 255949 263147 255984 263175
rect 255824 263113 255984 263147
rect 255824 263085 255859 263113
rect 255887 263085 255921 263113
rect 255949 263085 255984 263113
rect 255824 263051 255984 263085
rect 255824 263023 255859 263051
rect 255887 263023 255921 263051
rect 255949 263023 255984 263051
rect 255824 262989 255984 263023
rect 255824 262961 255859 262989
rect 255887 262961 255921 262989
rect 255949 262961 255984 262989
rect 255824 262944 255984 262961
rect 271184 263175 271344 263192
rect 271184 263147 271219 263175
rect 271247 263147 271281 263175
rect 271309 263147 271344 263175
rect 271184 263113 271344 263147
rect 271184 263085 271219 263113
rect 271247 263085 271281 263113
rect 271309 263085 271344 263113
rect 271184 263051 271344 263085
rect 271184 263023 271219 263051
rect 271247 263023 271281 263051
rect 271309 263023 271344 263051
rect 271184 262989 271344 263023
rect 271184 262961 271219 262989
rect 271247 262961 271281 262989
rect 271309 262961 271344 262989
rect 271184 262944 271344 262961
rect 279189 263175 279499 271961
rect 279189 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 279499 263175
rect 279189 263113 279499 263147
rect 279189 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 279499 263113
rect 279189 263051 279499 263085
rect 279189 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 279499 263051
rect 279189 262989 279499 263023
rect 279189 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 279499 262989
rect 98686 166553 98714 166558
rect 98742 260218 98770 260223
rect 98630 81881 98658 81886
rect 98686 164122 98714 164127
rect 96729 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 97039 77175
rect 96729 77113 97039 77147
rect 96729 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 97039 77113
rect 96729 77051 97039 77085
rect 96729 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 97039 77051
rect 96729 76989 97039 77023
rect 96729 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 97039 76989
rect 96729 68175 97039 76961
rect 96729 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 97039 68175
rect 96729 68113 97039 68147
rect 96729 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 97039 68113
rect 96729 68051 97039 68085
rect 96729 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 97039 68051
rect 96729 67989 97039 68023
rect 96729 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 97039 67989
rect 96729 59175 97039 67961
rect 98686 60746 98714 164094
rect 98742 152474 98770 260190
rect 109904 257175 110064 257192
rect 109904 257147 109939 257175
rect 109967 257147 110001 257175
rect 110029 257147 110064 257175
rect 109904 257113 110064 257147
rect 109904 257085 109939 257113
rect 109967 257085 110001 257113
rect 110029 257085 110064 257113
rect 109904 257051 110064 257085
rect 109904 257023 109939 257051
rect 109967 257023 110001 257051
rect 110029 257023 110064 257051
rect 109904 256989 110064 257023
rect 109904 256961 109939 256989
rect 109967 256961 110001 256989
rect 110029 256961 110064 256989
rect 109904 256944 110064 256961
rect 125264 257175 125424 257192
rect 125264 257147 125299 257175
rect 125327 257147 125361 257175
rect 125389 257147 125424 257175
rect 125264 257113 125424 257147
rect 125264 257085 125299 257113
rect 125327 257085 125361 257113
rect 125389 257085 125424 257113
rect 125264 257051 125424 257085
rect 125264 257023 125299 257051
rect 125327 257023 125361 257051
rect 125389 257023 125424 257051
rect 125264 256989 125424 257023
rect 125264 256961 125299 256989
rect 125327 256961 125361 256989
rect 125389 256961 125424 256989
rect 125264 256944 125424 256961
rect 140624 257175 140784 257192
rect 140624 257147 140659 257175
rect 140687 257147 140721 257175
rect 140749 257147 140784 257175
rect 140624 257113 140784 257147
rect 140624 257085 140659 257113
rect 140687 257085 140721 257113
rect 140749 257085 140784 257113
rect 140624 257051 140784 257085
rect 140624 257023 140659 257051
rect 140687 257023 140721 257051
rect 140749 257023 140784 257051
rect 140624 256989 140784 257023
rect 140624 256961 140659 256989
rect 140687 256961 140721 256989
rect 140749 256961 140784 256989
rect 140624 256944 140784 256961
rect 155984 257175 156144 257192
rect 155984 257147 156019 257175
rect 156047 257147 156081 257175
rect 156109 257147 156144 257175
rect 155984 257113 156144 257147
rect 155984 257085 156019 257113
rect 156047 257085 156081 257113
rect 156109 257085 156144 257113
rect 155984 257051 156144 257085
rect 155984 257023 156019 257051
rect 156047 257023 156081 257051
rect 156109 257023 156144 257051
rect 155984 256989 156144 257023
rect 155984 256961 156019 256989
rect 156047 256961 156081 256989
rect 156109 256961 156144 256989
rect 155984 256944 156144 256961
rect 171344 257175 171504 257192
rect 171344 257147 171379 257175
rect 171407 257147 171441 257175
rect 171469 257147 171504 257175
rect 171344 257113 171504 257147
rect 171344 257085 171379 257113
rect 171407 257085 171441 257113
rect 171469 257085 171504 257113
rect 171344 257051 171504 257085
rect 171344 257023 171379 257051
rect 171407 257023 171441 257051
rect 171469 257023 171504 257051
rect 171344 256989 171504 257023
rect 171344 256961 171379 256989
rect 171407 256961 171441 256989
rect 171469 256961 171504 256989
rect 171344 256944 171504 256961
rect 186704 257175 186864 257192
rect 186704 257147 186739 257175
rect 186767 257147 186801 257175
rect 186829 257147 186864 257175
rect 186704 257113 186864 257147
rect 186704 257085 186739 257113
rect 186767 257085 186801 257113
rect 186829 257085 186864 257113
rect 186704 257051 186864 257085
rect 186704 257023 186739 257051
rect 186767 257023 186801 257051
rect 186829 257023 186864 257051
rect 186704 256989 186864 257023
rect 186704 256961 186739 256989
rect 186767 256961 186801 256989
rect 186829 256961 186864 256989
rect 186704 256944 186864 256961
rect 202064 257175 202224 257192
rect 202064 257147 202099 257175
rect 202127 257147 202161 257175
rect 202189 257147 202224 257175
rect 202064 257113 202224 257147
rect 202064 257085 202099 257113
rect 202127 257085 202161 257113
rect 202189 257085 202224 257113
rect 202064 257051 202224 257085
rect 202064 257023 202099 257051
rect 202127 257023 202161 257051
rect 202189 257023 202224 257051
rect 202064 256989 202224 257023
rect 202064 256961 202099 256989
rect 202127 256961 202161 256989
rect 202189 256961 202224 256989
rect 202064 256944 202224 256961
rect 217424 257175 217584 257192
rect 217424 257147 217459 257175
rect 217487 257147 217521 257175
rect 217549 257147 217584 257175
rect 217424 257113 217584 257147
rect 217424 257085 217459 257113
rect 217487 257085 217521 257113
rect 217549 257085 217584 257113
rect 217424 257051 217584 257085
rect 217424 257023 217459 257051
rect 217487 257023 217521 257051
rect 217549 257023 217584 257051
rect 217424 256989 217584 257023
rect 217424 256961 217459 256989
rect 217487 256961 217521 256989
rect 217549 256961 217584 256989
rect 217424 256944 217584 256961
rect 232784 257175 232944 257192
rect 232784 257147 232819 257175
rect 232847 257147 232881 257175
rect 232909 257147 232944 257175
rect 232784 257113 232944 257147
rect 232784 257085 232819 257113
rect 232847 257085 232881 257113
rect 232909 257085 232944 257113
rect 232784 257051 232944 257085
rect 232784 257023 232819 257051
rect 232847 257023 232881 257051
rect 232909 257023 232944 257051
rect 232784 256989 232944 257023
rect 232784 256961 232819 256989
rect 232847 256961 232881 256989
rect 232909 256961 232944 256989
rect 232784 256944 232944 256961
rect 248144 257175 248304 257192
rect 248144 257147 248179 257175
rect 248207 257147 248241 257175
rect 248269 257147 248304 257175
rect 248144 257113 248304 257147
rect 248144 257085 248179 257113
rect 248207 257085 248241 257113
rect 248269 257085 248304 257113
rect 248144 257051 248304 257085
rect 248144 257023 248179 257051
rect 248207 257023 248241 257051
rect 248269 257023 248304 257051
rect 248144 256989 248304 257023
rect 248144 256961 248179 256989
rect 248207 256961 248241 256989
rect 248269 256961 248304 256989
rect 248144 256944 248304 256961
rect 263504 257175 263664 257192
rect 263504 257147 263539 257175
rect 263567 257147 263601 257175
rect 263629 257147 263664 257175
rect 263504 257113 263664 257147
rect 263504 257085 263539 257113
rect 263567 257085 263601 257113
rect 263629 257085 263664 257113
rect 263504 257051 263664 257085
rect 263504 257023 263539 257051
rect 263567 257023 263601 257051
rect 263629 257023 263664 257051
rect 263504 256989 263664 257023
rect 263504 256961 263539 256989
rect 263567 256961 263601 256989
rect 263629 256961 263664 256989
rect 263504 256944 263664 256961
rect 278864 257175 279024 257192
rect 278864 257147 278899 257175
rect 278927 257147 278961 257175
rect 278989 257147 279024 257175
rect 278864 257113 279024 257147
rect 278864 257085 278899 257113
rect 278927 257085 278961 257113
rect 278989 257085 279024 257113
rect 278864 257051 279024 257085
rect 278864 257023 278899 257051
rect 278927 257023 278961 257051
rect 278989 257023 279024 257051
rect 278864 256989 279024 257023
rect 278864 256961 278899 256989
rect 278927 256961 278961 256989
rect 278989 256961 279024 256989
rect 278864 256944 279024 256961
rect 102224 254175 102384 254192
rect 102224 254147 102259 254175
rect 102287 254147 102321 254175
rect 102349 254147 102384 254175
rect 102224 254113 102384 254147
rect 102224 254085 102259 254113
rect 102287 254085 102321 254113
rect 102349 254085 102384 254113
rect 102224 254051 102384 254085
rect 102224 254023 102259 254051
rect 102287 254023 102321 254051
rect 102349 254023 102384 254051
rect 102224 253989 102384 254023
rect 102224 253961 102259 253989
rect 102287 253961 102321 253989
rect 102349 253961 102384 253989
rect 102224 253944 102384 253961
rect 117584 254175 117744 254192
rect 117584 254147 117619 254175
rect 117647 254147 117681 254175
rect 117709 254147 117744 254175
rect 117584 254113 117744 254147
rect 117584 254085 117619 254113
rect 117647 254085 117681 254113
rect 117709 254085 117744 254113
rect 117584 254051 117744 254085
rect 117584 254023 117619 254051
rect 117647 254023 117681 254051
rect 117709 254023 117744 254051
rect 117584 253989 117744 254023
rect 117584 253961 117619 253989
rect 117647 253961 117681 253989
rect 117709 253961 117744 253989
rect 117584 253944 117744 253961
rect 132944 254175 133104 254192
rect 132944 254147 132979 254175
rect 133007 254147 133041 254175
rect 133069 254147 133104 254175
rect 132944 254113 133104 254147
rect 132944 254085 132979 254113
rect 133007 254085 133041 254113
rect 133069 254085 133104 254113
rect 132944 254051 133104 254085
rect 132944 254023 132979 254051
rect 133007 254023 133041 254051
rect 133069 254023 133104 254051
rect 132944 253989 133104 254023
rect 132944 253961 132979 253989
rect 133007 253961 133041 253989
rect 133069 253961 133104 253989
rect 132944 253944 133104 253961
rect 148304 254175 148464 254192
rect 148304 254147 148339 254175
rect 148367 254147 148401 254175
rect 148429 254147 148464 254175
rect 148304 254113 148464 254147
rect 148304 254085 148339 254113
rect 148367 254085 148401 254113
rect 148429 254085 148464 254113
rect 148304 254051 148464 254085
rect 148304 254023 148339 254051
rect 148367 254023 148401 254051
rect 148429 254023 148464 254051
rect 148304 253989 148464 254023
rect 148304 253961 148339 253989
rect 148367 253961 148401 253989
rect 148429 253961 148464 253989
rect 148304 253944 148464 253961
rect 163664 254175 163824 254192
rect 163664 254147 163699 254175
rect 163727 254147 163761 254175
rect 163789 254147 163824 254175
rect 163664 254113 163824 254147
rect 163664 254085 163699 254113
rect 163727 254085 163761 254113
rect 163789 254085 163824 254113
rect 163664 254051 163824 254085
rect 163664 254023 163699 254051
rect 163727 254023 163761 254051
rect 163789 254023 163824 254051
rect 163664 253989 163824 254023
rect 163664 253961 163699 253989
rect 163727 253961 163761 253989
rect 163789 253961 163824 253989
rect 163664 253944 163824 253961
rect 179024 254175 179184 254192
rect 179024 254147 179059 254175
rect 179087 254147 179121 254175
rect 179149 254147 179184 254175
rect 179024 254113 179184 254147
rect 179024 254085 179059 254113
rect 179087 254085 179121 254113
rect 179149 254085 179184 254113
rect 179024 254051 179184 254085
rect 179024 254023 179059 254051
rect 179087 254023 179121 254051
rect 179149 254023 179184 254051
rect 179024 253989 179184 254023
rect 179024 253961 179059 253989
rect 179087 253961 179121 253989
rect 179149 253961 179184 253989
rect 179024 253944 179184 253961
rect 194384 254175 194544 254192
rect 194384 254147 194419 254175
rect 194447 254147 194481 254175
rect 194509 254147 194544 254175
rect 194384 254113 194544 254147
rect 194384 254085 194419 254113
rect 194447 254085 194481 254113
rect 194509 254085 194544 254113
rect 194384 254051 194544 254085
rect 194384 254023 194419 254051
rect 194447 254023 194481 254051
rect 194509 254023 194544 254051
rect 194384 253989 194544 254023
rect 194384 253961 194419 253989
rect 194447 253961 194481 253989
rect 194509 253961 194544 253989
rect 194384 253944 194544 253961
rect 209744 254175 209904 254192
rect 209744 254147 209779 254175
rect 209807 254147 209841 254175
rect 209869 254147 209904 254175
rect 209744 254113 209904 254147
rect 209744 254085 209779 254113
rect 209807 254085 209841 254113
rect 209869 254085 209904 254113
rect 209744 254051 209904 254085
rect 209744 254023 209779 254051
rect 209807 254023 209841 254051
rect 209869 254023 209904 254051
rect 209744 253989 209904 254023
rect 209744 253961 209779 253989
rect 209807 253961 209841 253989
rect 209869 253961 209904 253989
rect 209744 253944 209904 253961
rect 225104 254175 225264 254192
rect 225104 254147 225139 254175
rect 225167 254147 225201 254175
rect 225229 254147 225264 254175
rect 225104 254113 225264 254147
rect 225104 254085 225139 254113
rect 225167 254085 225201 254113
rect 225229 254085 225264 254113
rect 225104 254051 225264 254085
rect 225104 254023 225139 254051
rect 225167 254023 225201 254051
rect 225229 254023 225264 254051
rect 225104 253989 225264 254023
rect 225104 253961 225139 253989
rect 225167 253961 225201 253989
rect 225229 253961 225264 253989
rect 225104 253944 225264 253961
rect 240464 254175 240624 254192
rect 240464 254147 240499 254175
rect 240527 254147 240561 254175
rect 240589 254147 240624 254175
rect 240464 254113 240624 254147
rect 240464 254085 240499 254113
rect 240527 254085 240561 254113
rect 240589 254085 240624 254113
rect 240464 254051 240624 254085
rect 240464 254023 240499 254051
rect 240527 254023 240561 254051
rect 240589 254023 240624 254051
rect 240464 253989 240624 254023
rect 240464 253961 240499 253989
rect 240527 253961 240561 253989
rect 240589 253961 240624 253989
rect 240464 253944 240624 253961
rect 255824 254175 255984 254192
rect 255824 254147 255859 254175
rect 255887 254147 255921 254175
rect 255949 254147 255984 254175
rect 255824 254113 255984 254147
rect 255824 254085 255859 254113
rect 255887 254085 255921 254113
rect 255949 254085 255984 254113
rect 255824 254051 255984 254085
rect 255824 254023 255859 254051
rect 255887 254023 255921 254051
rect 255949 254023 255984 254051
rect 255824 253989 255984 254023
rect 255824 253961 255859 253989
rect 255887 253961 255921 253989
rect 255949 253961 255984 253989
rect 255824 253944 255984 253961
rect 271184 254175 271344 254192
rect 271184 254147 271219 254175
rect 271247 254147 271281 254175
rect 271309 254147 271344 254175
rect 271184 254113 271344 254147
rect 271184 254085 271219 254113
rect 271247 254085 271281 254113
rect 271309 254085 271344 254113
rect 271184 254051 271344 254085
rect 271184 254023 271219 254051
rect 271247 254023 271281 254051
rect 271309 254023 271344 254051
rect 271184 253989 271344 254023
rect 271184 253961 271219 253989
rect 271247 253961 271281 253989
rect 271309 253961 271344 253989
rect 271184 253944 271344 253961
rect 279189 254175 279499 262961
rect 279189 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 279499 254175
rect 279189 254113 279499 254147
rect 279189 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 279499 254113
rect 279189 254051 279499 254085
rect 279189 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 279499 254051
rect 279189 253989 279499 254023
rect 279189 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 279499 253989
rect 98854 252826 98882 252831
rect 98742 152441 98770 152446
rect 98798 230650 98826 230655
rect 98686 60713 98714 60718
rect 98742 149338 98770 149343
rect 96729 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 97039 59175
rect 96729 59113 97039 59147
rect 96729 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 97039 59113
rect 96729 59051 97039 59085
rect 96729 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 97039 59051
rect 96729 58989 97039 59023
rect 96729 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 97039 58989
rect 96729 50175 97039 58961
rect 96729 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 97039 50175
rect 96729 50113 97039 50147
rect 96729 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 97039 50113
rect 96729 50051 97039 50085
rect 96729 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 97039 50051
rect 96729 49989 97039 50023
rect 96729 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 97039 49989
rect 96729 41175 97039 49961
rect 98742 46634 98770 149310
rect 98798 124250 98826 230622
rect 98854 145418 98882 252798
rect 109904 248175 110064 248192
rect 109904 248147 109939 248175
rect 109967 248147 110001 248175
rect 110029 248147 110064 248175
rect 109904 248113 110064 248147
rect 109904 248085 109939 248113
rect 109967 248085 110001 248113
rect 110029 248085 110064 248113
rect 109904 248051 110064 248085
rect 109904 248023 109939 248051
rect 109967 248023 110001 248051
rect 110029 248023 110064 248051
rect 109904 247989 110064 248023
rect 109904 247961 109939 247989
rect 109967 247961 110001 247989
rect 110029 247961 110064 247989
rect 109904 247944 110064 247961
rect 125264 248175 125424 248192
rect 125264 248147 125299 248175
rect 125327 248147 125361 248175
rect 125389 248147 125424 248175
rect 125264 248113 125424 248147
rect 125264 248085 125299 248113
rect 125327 248085 125361 248113
rect 125389 248085 125424 248113
rect 125264 248051 125424 248085
rect 125264 248023 125299 248051
rect 125327 248023 125361 248051
rect 125389 248023 125424 248051
rect 125264 247989 125424 248023
rect 125264 247961 125299 247989
rect 125327 247961 125361 247989
rect 125389 247961 125424 247989
rect 125264 247944 125424 247961
rect 140624 248175 140784 248192
rect 140624 248147 140659 248175
rect 140687 248147 140721 248175
rect 140749 248147 140784 248175
rect 140624 248113 140784 248147
rect 140624 248085 140659 248113
rect 140687 248085 140721 248113
rect 140749 248085 140784 248113
rect 140624 248051 140784 248085
rect 140624 248023 140659 248051
rect 140687 248023 140721 248051
rect 140749 248023 140784 248051
rect 140624 247989 140784 248023
rect 140624 247961 140659 247989
rect 140687 247961 140721 247989
rect 140749 247961 140784 247989
rect 140624 247944 140784 247961
rect 155984 248175 156144 248192
rect 155984 248147 156019 248175
rect 156047 248147 156081 248175
rect 156109 248147 156144 248175
rect 155984 248113 156144 248147
rect 155984 248085 156019 248113
rect 156047 248085 156081 248113
rect 156109 248085 156144 248113
rect 155984 248051 156144 248085
rect 155984 248023 156019 248051
rect 156047 248023 156081 248051
rect 156109 248023 156144 248051
rect 155984 247989 156144 248023
rect 155984 247961 156019 247989
rect 156047 247961 156081 247989
rect 156109 247961 156144 247989
rect 155984 247944 156144 247961
rect 171344 248175 171504 248192
rect 171344 248147 171379 248175
rect 171407 248147 171441 248175
rect 171469 248147 171504 248175
rect 171344 248113 171504 248147
rect 171344 248085 171379 248113
rect 171407 248085 171441 248113
rect 171469 248085 171504 248113
rect 171344 248051 171504 248085
rect 171344 248023 171379 248051
rect 171407 248023 171441 248051
rect 171469 248023 171504 248051
rect 171344 247989 171504 248023
rect 171344 247961 171379 247989
rect 171407 247961 171441 247989
rect 171469 247961 171504 247989
rect 171344 247944 171504 247961
rect 186704 248175 186864 248192
rect 186704 248147 186739 248175
rect 186767 248147 186801 248175
rect 186829 248147 186864 248175
rect 186704 248113 186864 248147
rect 186704 248085 186739 248113
rect 186767 248085 186801 248113
rect 186829 248085 186864 248113
rect 186704 248051 186864 248085
rect 186704 248023 186739 248051
rect 186767 248023 186801 248051
rect 186829 248023 186864 248051
rect 186704 247989 186864 248023
rect 186704 247961 186739 247989
rect 186767 247961 186801 247989
rect 186829 247961 186864 247989
rect 186704 247944 186864 247961
rect 202064 248175 202224 248192
rect 202064 248147 202099 248175
rect 202127 248147 202161 248175
rect 202189 248147 202224 248175
rect 202064 248113 202224 248147
rect 202064 248085 202099 248113
rect 202127 248085 202161 248113
rect 202189 248085 202224 248113
rect 202064 248051 202224 248085
rect 202064 248023 202099 248051
rect 202127 248023 202161 248051
rect 202189 248023 202224 248051
rect 202064 247989 202224 248023
rect 202064 247961 202099 247989
rect 202127 247961 202161 247989
rect 202189 247961 202224 247989
rect 202064 247944 202224 247961
rect 217424 248175 217584 248192
rect 217424 248147 217459 248175
rect 217487 248147 217521 248175
rect 217549 248147 217584 248175
rect 217424 248113 217584 248147
rect 217424 248085 217459 248113
rect 217487 248085 217521 248113
rect 217549 248085 217584 248113
rect 217424 248051 217584 248085
rect 217424 248023 217459 248051
rect 217487 248023 217521 248051
rect 217549 248023 217584 248051
rect 217424 247989 217584 248023
rect 217424 247961 217459 247989
rect 217487 247961 217521 247989
rect 217549 247961 217584 247989
rect 217424 247944 217584 247961
rect 232784 248175 232944 248192
rect 232784 248147 232819 248175
rect 232847 248147 232881 248175
rect 232909 248147 232944 248175
rect 232784 248113 232944 248147
rect 232784 248085 232819 248113
rect 232847 248085 232881 248113
rect 232909 248085 232944 248113
rect 232784 248051 232944 248085
rect 232784 248023 232819 248051
rect 232847 248023 232881 248051
rect 232909 248023 232944 248051
rect 232784 247989 232944 248023
rect 232784 247961 232819 247989
rect 232847 247961 232881 247989
rect 232909 247961 232944 247989
rect 232784 247944 232944 247961
rect 248144 248175 248304 248192
rect 248144 248147 248179 248175
rect 248207 248147 248241 248175
rect 248269 248147 248304 248175
rect 248144 248113 248304 248147
rect 248144 248085 248179 248113
rect 248207 248085 248241 248113
rect 248269 248085 248304 248113
rect 248144 248051 248304 248085
rect 248144 248023 248179 248051
rect 248207 248023 248241 248051
rect 248269 248023 248304 248051
rect 248144 247989 248304 248023
rect 248144 247961 248179 247989
rect 248207 247961 248241 247989
rect 248269 247961 248304 247989
rect 248144 247944 248304 247961
rect 263504 248175 263664 248192
rect 263504 248147 263539 248175
rect 263567 248147 263601 248175
rect 263629 248147 263664 248175
rect 263504 248113 263664 248147
rect 263504 248085 263539 248113
rect 263567 248085 263601 248113
rect 263629 248085 263664 248113
rect 263504 248051 263664 248085
rect 263504 248023 263539 248051
rect 263567 248023 263601 248051
rect 263629 248023 263664 248051
rect 263504 247989 263664 248023
rect 263504 247961 263539 247989
rect 263567 247961 263601 247989
rect 263629 247961 263664 247989
rect 263504 247944 263664 247961
rect 278864 248175 279024 248192
rect 278864 248147 278899 248175
rect 278927 248147 278961 248175
rect 278989 248147 279024 248175
rect 278864 248113 279024 248147
rect 278864 248085 278899 248113
rect 278927 248085 278961 248113
rect 278989 248085 279024 248113
rect 278864 248051 279024 248085
rect 278864 248023 278899 248051
rect 278927 248023 278961 248051
rect 278989 248023 279024 248051
rect 278864 247989 279024 248023
rect 278864 247961 278899 247989
rect 278927 247961 278961 247989
rect 278989 247961 279024 247989
rect 278864 247944 279024 247961
rect 102224 245175 102384 245192
rect 102224 245147 102259 245175
rect 102287 245147 102321 245175
rect 102349 245147 102384 245175
rect 102224 245113 102384 245147
rect 102224 245085 102259 245113
rect 102287 245085 102321 245113
rect 102349 245085 102384 245113
rect 102224 245051 102384 245085
rect 102224 245023 102259 245051
rect 102287 245023 102321 245051
rect 102349 245023 102384 245051
rect 102224 244989 102384 245023
rect 102224 244961 102259 244989
rect 102287 244961 102321 244989
rect 102349 244961 102384 244989
rect 102224 244944 102384 244961
rect 117584 245175 117744 245192
rect 117584 245147 117619 245175
rect 117647 245147 117681 245175
rect 117709 245147 117744 245175
rect 117584 245113 117744 245147
rect 117584 245085 117619 245113
rect 117647 245085 117681 245113
rect 117709 245085 117744 245113
rect 117584 245051 117744 245085
rect 117584 245023 117619 245051
rect 117647 245023 117681 245051
rect 117709 245023 117744 245051
rect 117584 244989 117744 245023
rect 117584 244961 117619 244989
rect 117647 244961 117681 244989
rect 117709 244961 117744 244989
rect 117584 244944 117744 244961
rect 132944 245175 133104 245192
rect 132944 245147 132979 245175
rect 133007 245147 133041 245175
rect 133069 245147 133104 245175
rect 132944 245113 133104 245147
rect 132944 245085 132979 245113
rect 133007 245085 133041 245113
rect 133069 245085 133104 245113
rect 132944 245051 133104 245085
rect 132944 245023 132979 245051
rect 133007 245023 133041 245051
rect 133069 245023 133104 245051
rect 132944 244989 133104 245023
rect 132944 244961 132979 244989
rect 133007 244961 133041 244989
rect 133069 244961 133104 244989
rect 132944 244944 133104 244961
rect 148304 245175 148464 245192
rect 148304 245147 148339 245175
rect 148367 245147 148401 245175
rect 148429 245147 148464 245175
rect 148304 245113 148464 245147
rect 148304 245085 148339 245113
rect 148367 245085 148401 245113
rect 148429 245085 148464 245113
rect 148304 245051 148464 245085
rect 148304 245023 148339 245051
rect 148367 245023 148401 245051
rect 148429 245023 148464 245051
rect 148304 244989 148464 245023
rect 148304 244961 148339 244989
rect 148367 244961 148401 244989
rect 148429 244961 148464 244989
rect 148304 244944 148464 244961
rect 163664 245175 163824 245192
rect 163664 245147 163699 245175
rect 163727 245147 163761 245175
rect 163789 245147 163824 245175
rect 163664 245113 163824 245147
rect 163664 245085 163699 245113
rect 163727 245085 163761 245113
rect 163789 245085 163824 245113
rect 163664 245051 163824 245085
rect 163664 245023 163699 245051
rect 163727 245023 163761 245051
rect 163789 245023 163824 245051
rect 163664 244989 163824 245023
rect 163664 244961 163699 244989
rect 163727 244961 163761 244989
rect 163789 244961 163824 244989
rect 163664 244944 163824 244961
rect 179024 245175 179184 245192
rect 179024 245147 179059 245175
rect 179087 245147 179121 245175
rect 179149 245147 179184 245175
rect 179024 245113 179184 245147
rect 179024 245085 179059 245113
rect 179087 245085 179121 245113
rect 179149 245085 179184 245113
rect 179024 245051 179184 245085
rect 179024 245023 179059 245051
rect 179087 245023 179121 245051
rect 179149 245023 179184 245051
rect 179024 244989 179184 245023
rect 179024 244961 179059 244989
rect 179087 244961 179121 244989
rect 179149 244961 179184 244989
rect 179024 244944 179184 244961
rect 194384 245175 194544 245192
rect 194384 245147 194419 245175
rect 194447 245147 194481 245175
rect 194509 245147 194544 245175
rect 194384 245113 194544 245147
rect 194384 245085 194419 245113
rect 194447 245085 194481 245113
rect 194509 245085 194544 245113
rect 194384 245051 194544 245085
rect 194384 245023 194419 245051
rect 194447 245023 194481 245051
rect 194509 245023 194544 245051
rect 194384 244989 194544 245023
rect 194384 244961 194419 244989
rect 194447 244961 194481 244989
rect 194509 244961 194544 244989
rect 194384 244944 194544 244961
rect 209744 245175 209904 245192
rect 209744 245147 209779 245175
rect 209807 245147 209841 245175
rect 209869 245147 209904 245175
rect 209744 245113 209904 245147
rect 209744 245085 209779 245113
rect 209807 245085 209841 245113
rect 209869 245085 209904 245113
rect 209744 245051 209904 245085
rect 209744 245023 209779 245051
rect 209807 245023 209841 245051
rect 209869 245023 209904 245051
rect 209744 244989 209904 245023
rect 209744 244961 209779 244989
rect 209807 244961 209841 244989
rect 209869 244961 209904 244989
rect 209744 244944 209904 244961
rect 225104 245175 225264 245192
rect 225104 245147 225139 245175
rect 225167 245147 225201 245175
rect 225229 245147 225264 245175
rect 225104 245113 225264 245147
rect 225104 245085 225139 245113
rect 225167 245085 225201 245113
rect 225229 245085 225264 245113
rect 225104 245051 225264 245085
rect 225104 245023 225139 245051
rect 225167 245023 225201 245051
rect 225229 245023 225264 245051
rect 225104 244989 225264 245023
rect 225104 244961 225139 244989
rect 225167 244961 225201 244989
rect 225229 244961 225264 244989
rect 225104 244944 225264 244961
rect 240464 245175 240624 245192
rect 240464 245147 240499 245175
rect 240527 245147 240561 245175
rect 240589 245147 240624 245175
rect 240464 245113 240624 245147
rect 240464 245085 240499 245113
rect 240527 245085 240561 245113
rect 240589 245085 240624 245113
rect 240464 245051 240624 245085
rect 240464 245023 240499 245051
rect 240527 245023 240561 245051
rect 240589 245023 240624 245051
rect 240464 244989 240624 245023
rect 240464 244961 240499 244989
rect 240527 244961 240561 244989
rect 240589 244961 240624 244989
rect 240464 244944 240624 244961
rect 255824 245175 255984 245192
rect 255824 245147 255859 245175
rect 255887 245147 255921 245175
rect 255949 245147 255984 245175
rect 255824 245113 255984 245147
rect 255824 245085 255859 245113
rect 255887 245085 255921 245113
rect 255949 245085 255984 245113
rect 255824 245051 255984 245085
rect 255824 245023 255859 245051
rect 255887 245023 255921 245051
rect 255949 245023 255984 245051
rect 255824 244989 255984 245023
rect 255824 244961 255859 244989
rect 255887 244961 255921 244989
rect 255949 244961 255984 244989
rect 255824 244944 255984 244961
rect 271184 245175 271344 245192
rect 271184 245147 271219 245175
rect 271247 245147 271281 245175
rect 271309 245147 271344 245175
rect 271184 245113 271344 245147
rect 271184 245085 271219 245113
rect 271247 245085 271281 245113
rect 271309 245085 271344 245113
rect 271184 245051 271344 245085
rect 271184 245023 271219 245051
rect 271247 245023 271281 245051
rect 271309 245023 271344 245051
rect 271184 244989 271344 245023
rect 271184 244961 271219 244989
rect 271247 244961 271281 244989
rect 271309 244961 271344 244989
rect 271184 244944 271344 244961
rect 279189 245175 279499 253961
rect 279189 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 279499 245175
rect 279189 245113 279499 245147
rect 279189 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 279499 245113
rect 279189 245051 279499 245085
rect 279189 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 279499 245051
rect 279189 244989 279499 245023
rect 279189 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 279499 244989
rect 109904 239175 110064 239192
rect 109904 239147 109939 239175
rect 109967 239147 110001 239175
rect 110029 239147 110064 239175
rect 109904 239113 110064 239147
rect 109904 239085 109939 239113
rect 109967 239085 110001 239113
rect 110029 239085 110064 239113
rect 109904 239051 110064 239085
rect 109904 239023 109939 239051
rect 109967 239023 110001 239051
rect 110029 239023 110064 239051
rect 109904 238989 110064 239023
rect 109904 238961 109939 238989
rect 109967 238961 110001 238989
rect 110029 238961 110064 238989
rect 109904 238944 110064 238961
rect 125264 239175 125424 239192
rect 125264 239147 125299 239175
rect 125327 239147 125361 239175
rect 125389 239147 125424 239175
rect 125264 239113 125424 239147
rect 125264 239085 125299 239113
rect 125327 239085 125361 239113
rect 125389 239085 125424 239113
rect 125264 239051 125424 239085
rect 125264 239023 125299 239051
rect 125327 239023 125361 239051
rect 125389 239023 125424 239051
rect 125264 238989 125424 239023
rect 125264 238961 125299 238989
rect 125327 238961 125361 238989
rect 125389 238961 125424 238989
rect 125264 238944 125424 238961
rect 140624 239175 140784 239192
rect 140624 239147 140659 239175
rect 140687 239147 140721 239175
rect 140749 239147 140784 239175
rect 140624 239113 140784 239147
rect 140624 239085 140659 239113
rect 140687 239085 140721 239113
rect 140749 239085 140784 239113
rect 140624 239051 140784 239085
rect 140624 239023 140659 239051
rect 140687 239023 140721 239051
rect 140749 239023 140784 239051
rect 140624 238989 140784 239023
rect 140624 238961 140659 238989
rect 140687 238961 140721 238989
rect 140749 238961 140784 238989
rect 140624 238944 140784 238961
rect 155984 239175 156144 239192
rect 155984 239147 156019 239175
rect 156047 239147 156081 239175
rect 156109 239147 156144 239175
rect 155984 239113 156144 239147
rect 155984 239085 156019 239113
rect 156047 239085 156081 239113
rect 156109 239085 156144 239113
rect 155984 239051 156144 239085
rect 155984 239023 156019 239051
rect 156047 239023 156081 239051
rect 156109 239023 156144 239051
rect 155984 238989 156144 239023
rect 155984 238961 156019 238989
rect 156047 238961 156081 238989
rect 156109 238961 156144 238989
rect 155984 238944 156144 238961
rect 171344 239175 171504 239192
rect 171344 239147 171379 239175
rect 171407 239147 171441 239175
rect 171469 239147 171504 239175
rect 171344 239113 171504 239147
rect 171344 239085 171379 239113
rect 171407 239085 171441 239113
rect 171469 239085 171504 239113
rect 171344 239051 171504 239085
rect 171344 239023 171379 239051
rect 171407 239023 171441 239051
rect 171469 239023 171504 239051
rect 171344 238989 171504 239023
rect 171344 238961 171379 238989
rect 171407 238961 171441 238989
rect 171469 238961 171504 238989
rect 171344 238944 171504 238961
rect 186704 239175 186864 239192
rect 186704 239147 186739 239175
rect 186767 239147 186801 239175
rect 186829 239147 186864 239175
rect 186704 239113 186864 239147
rect 186704 239085 186739 239113
rect 186767 239085 186801 239113
rect 186829 239085 186864 239113
rect 186704 239051 186864 239085
rect 186704 239023 186739 239051
rect 186767 239023 186801 239051
rect 186829 239023 186864 239051
rect 186704 238989 186864 239023
rect 186704 238961 186739 238989
rect 186767 238961 186801 238989
rect 186829 238961 186864 238989
rect 186704 238944 186864 238961
rect 202064 239175 202224 239192
rect 202064 239147 202099 239175
rect 202127 239147 202161 239175
rect 202189 239147 202224 239175
rect 202064 239113 202224 239147
rect 202064 239085 202099 239113
rect 202127 239085 202161 239113
rect 202189 239085 202224 239113
rect 202064 239051 202224 239085
rect 202064 239023 202099 239051
rect 202127 239023 202161 239051
rect 202189 239023 202224 239051
rect 202064 238989 202224 239023
rect 202064 238961 202099 238989
rect 202127 238961 202161 238989
rect 202189 238961 202224 238989
rect 202064 238944 202224 238961
rect 217424 239175 217584 239192
rect 217424 239147 217459 239175
rect 217487 239147 217521 239175
rect 217549 239147 217584 239175
rect 217424 239113 217584 239147
rect 217424 239085 217459 239113
rect 217487 239085 217521 239113
rect 217549 239085 217584 239113
rect 217424 239051 217584 239085
rect 217424 239023 217459 239051
rect 217487 239023 217521 239051
rect 217549 239023 217584 239051
rect 217424 238989 217584 239023
rect 217424 238961 217459 238989
rect 217487 238961 217521 238989
rect 217549 238961 217584 238989
rect 217424 238944 217584 238961
rect 232784 239175 232944 239192
rect 232784 239147 232819 239175
rect 232847 239147 232881 239175
rect 232909 239147 232944 239175
rect 232784 239113 232944 239147
rect 232784 239085 232819 239113
rect 232847 239085 232881 239113
rect 232909 239085 232944 239113
rect 232784 239051 232944 239085
rect 232784 239023 232819 239051
rect 232847 239023 232881 239051
rect 232909 239023 232944 239051
rect 232784 238989 232944 239023
rect 232784 238961 232819 238989
rect 232847 238961 232881 238989
rect 232909 238961 232944 238989
rect 232784 238944 232944 238961
rect 248144 239175 248304 239192
rect 248144 239147 248179 239175
rect 248207 239147 248241 239175
rect 248269 239147 248304 239175
rect 248144 239113 248304 239147
rect 248144 239085 248179 239113
rect 248207 239085 248241 239113
rect 248269 239085 248304 239113
rect 248144 239051 248304 239085
rect 248144 239023 248179 239051
rect 248207 239023 248241 239051
rect 248269 239023 248304 239051
rect 248144 238989 248304 239023
rect 248144 238961 248179 238989
rect 248207 238961 248241 238989
rect 248269 238961 248304 238989
rect 248144 238944 248304 238961
rect 263504 239175 263664 239192
rect 263504 239147 263539 239175
rect 263567 239147 263601 239175
rect 263629 239147 263664 239175
rect 263504 239113 263664 239147
rect 263504 239085 263539 239113
rect 263567 239085 263601 239113
rect 263629 239085 263664 239113
rect 263504 239051 263664 239085
rect 263504 239023 263539 239051
rect 263567 239023 263601 239051
rect 263629 239023 263664 239051
rect 263504 238989 263664 239023
rect 263504 238961 263539 238989
rect 263567 238961 263601 238989
rect 263629 238961 263664 238989
rect 263504 238944 263664 238961
rect 278864 239175 279024 239192
rect 278864 239147 278899 239175
rect 278927 239147 278961 239175
rect 278989 239147 279024 239175
rect 278864 239113 279024 239147
rect 278864 239085 278899 239113
rect 278927 239085 278961 239113
rect 278989 239085 279024 239113
rect 278864 239051 279024 239085
rect 278864 239023 278899 239051
rect 278927 239023 278961 239051
rect 278989 239023 279024 239051
rect 278864 238989 279024 239023
rect 278864 238961 278899 238989
rect 278927 238961 278961 238989
rect 278989 238961 279024 238989
rect 278864 238944 279024 238961
rect 102224 236175 102384 236192
rect 102224 236147 102259 236175
rect 102287 236147 102321 236175
rect 102349 236147 102384 236175
rect 102224 236113 102384 236147
rect 102224 236085 102259 236113
rect 102287 236085 102321 236113
rect 102349 236085 102384 236113
rect 102224 236051 102384 236085
rect 102224 236023 102259 236051
rect 102287 236023 102321 236051
rect 102349 236023 102384 236051
rect 102224 235989 102384 236023
rect 102224 235961 102259 235989
rect 102287 235961 102321 235989
rect 102349 235961 102384 235989
rect 102224 235944 102384 235961
rect 117584 236175 117744 236192
rect 117584 236147 117619 236175
rect 117647 236147 117681 236175
rect 117709 236147 117744 236175
rect 117584 236113 117744 236147
rect 117584 236085 117619 236113
rect 117647 236085 117681 236113
rect 117709 236085 117744 236113
rect 117584 236051 117744 236085
rect 117584 236023 117619 236051
rect 117647 236023 117681 236051
rect 117709 236023 117744 236051
rect 117584 235989 117744 236023
rect 117584 235961 117619 235989
rect 117647 235961 117681 235989
rect 117709 235961 117744 235989
rect 117584 235944 117744 235961
rect 132944 236175 133104 236192
rect 132944 236147 132979 236175
rect 133007 236147 133041 236175
rect 133069 236147 133104 236175
rect 132944 236113 133104 236147
rect 132944 236085 132979 236113
rect 133007 236085 133041 236113
rect 133069 236085 133104 236113
rect 132944 236051 133104 236085
rect 132944 236023 132979 236051
rect 133007 236023 133041 236051
rect 133069 236023 133104 236051
rect 132944 235989 133104 236023
rect 132944 235961 132979 235989
rect 133007 235961 133041 235989
rect 133069 235961 133104 235989
rect 132944 235944 133104 235961
rect 148304 236175 148464 236192
rect 148304 236147 148339 236175
rect 148367 236147 148401 236175
rect 148429 236147 148464 236175
rect 148304 236113 148464 236147
rect 148304 236085 148339 236113
rect 148367 236085 148401 236113
rect 148429 236085 148464 236113
rect 148304 236051 148464 236085
rect 148304 236023 148339 236051
rect 148367 236023 148401 236051
rect 148429 236023 148464 236051
rect 148304 235989 148464 236023
rect 148304 235961 148339 235989
rect 148367 235961 148401 235989
rect 148429 235961 148464 235989
rect 148304 235944 148464 235961
rect 163664 236175 163824 236192
rect 163664 236147 163699 236175
rect 163727 236147 163761 236175
rect 163789 236147 163824 236175
rect 163664 236113 163824 236147
rect 163664 236085 163699 236113
rect 163727 236085 163761 236113
rect 163789 236085 163824 236113
rect 163664 236051 163824 236085
rect 163664 236023 163699 236051
rect 163727 236023 163761 236051
rect 163789 236023 163824 236051
rect 163664 235989 163824 236023
rect 163664 235961 163699 235989
rect 163727 235961 163761 235989
rect 163789 235961 163824 235989
rect 163664 235944 163824 235961
rect 179024 236175 179184 236192
rect 179024 236147 179059 236175
rect 179087 236147 179121 236175
rect 179149 236147 179184 236175
rect 179024 236113 179184 236147
rect 179024 236085 179059 236113
rect 179087 236085 179121 236113
rect 179149 236085 179184 236113
rect 179024 236051 179184 236085
rect 179024 236023 179059 236051
rect 179087 236023 179121 236051
rect 179149 236023 179184 236051
rect 179024 235989 179184 236023
rect 179024 235961 179059 235989
rect 179087 235961 179121 235989
rect 179149 235961 179184 235989
rect 179024 235944 179184 235961
rect 194384 236175 194544 236192
rect 194384 236147 194419 236175
rect 194447 236147 194481 236175
rect 194509 236147 194544 236175
rect 194384 236113 194544 236147
rect 194384 236085 194419 236113
rect 194447 236085 194481 236113
rect 194509 236085 194544 236113
rect 194384 236051 194544 236085
rect 194384 236023 194419 236051
rect 194447 236023 194481 236051
rect 194509 236023 194544 236051
rect 194384 235989 194544 236023
rect 194384 235961 194419 235989
rect 194447 235961 194481 235989
rect 194509 235961 194544 235989
rect 194384 235944 194544 235961
rect 209744 236175 209904 236192
rect 209744 236147 209779 236175
rect 209807 236147 209841 236175
rect 209869 236147 209904 236175
rect 209744 236113 209904 236147
rect 209744 236085 209779 236113
rect 209807 236085 209841 236113
rect 209869 236085 209904 236113
rect 209744 236051 209904 236085
rect 209744 236023 209779 236051
rect 209807 236023 209841 236051
rect 209869 236023 209904 236051
rect 209744 235989 209904 236023
rect 209744 235961 209779 235989
rect 209807 235961 209841 235989
rect 209869 235961 209904 235989
rect 209744 235944 209904 235961
rect 225104 236175 225264 236192
rect 225104 236147 225139 236175
rect 225167 236147 225201 236175
rect 225229 236147 225264 236175
rect 225104 236113 225264 236147
rect 225104 236085 225139 236113
rect 225167 236085 225201 236113
rect 225229 236085 225264 236113
rect 225104 236051 225264 236085
rect 225104 236023 225139 236051
rect 225167 236023 225201 236051
rect 225229 236023 225264 236051
rect 225104 235989 225264 236023
rect 225104 235961 225139 235989
rect 225167 235961 225201 235989
rect 225229 235961 225264 235989
rect 225104 235944 225264 235961
rect 240464 236175 240624 236192
rect 240464 236147 240499 236175
rect 240527 236147 240561 236175
rect 240589 236147 240624 236175
rect 240464 236113 240624 236147
rect 240464 236085 240499 236113
rect 240527 236085 240561 236113
rect 240589 236085 240624 236113
rect 240464 236051 240624 236085
rect 240464 236023 240499 236051
rect 240527 236023 240561 236051
rect 240589 236023 240624 236051
rect 240464 235989 240624 236023
rect 240464 235961 240499 235989
rect 240527 235961 240561 235989
rect 240589 235961 240624 235989
rect 240464 235944 240624 235961
rect 255824 236175 255984 236192
rect 255824 236147 255859 236175
rect 255887 236147 255921 236175
rect 255949 236147 255984 236175
rect 255824 236113 255984 236147
rect 255824 236085 255859 236113
rect 255887 236085 255921 236113
rect 255949 236085 255984 236113
rect 255824 236051 255984 236085
rect 255824 236023 255859 236051
rect 255887 236023 255921 236051
rect 255949 236023 255984 236051
rect 255824 235989 255984 236023
rect 255824 235961 255859 235989
rect 255887 235961 255921 235989
rect 255949 235961 255984 235989
rect 255824 235944 255984 235961
rect 271184 236175 271344 236192
rect 271184 236147 271219 236175
rect 271247 236147 271281 236175
rect 271309 236147 271344 236175
rect 271184 236113 271344 236147
rect 271184 236085 271219 236113
rect 271247 236085 271281 236113
rect 271309 236085 271344 236113
rect 271184 236051 271344 236085
rect 271184 236023 271219 236051
rect 271247 236023 271281 236051
rect 271309 236023 271344 236051
rect 271184 235989 271344 236023
rect 271184 235961 271219 235989
rect 271247 235961 271281 235989
rect 271309 235961 271344 235989
rect 271184 235944 271344 235961
rect 279189 236175 279499 244961
rect 279189 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 279499 236175
rect 279189 236113 279499 236147
rect 279189 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 279499 236113
rect 279189 236051 279499 236085
rect 279189 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 279499 236051
rect 279189 235989 279499 236023
rect 279189 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 279499 235989
rect 109904 230175 110064 230192
rect 109904 230147 109939 230175
rect 109967 230147 110001 230175
rect 110029 230147 110064 230175
rect 109904 230113 110064 230147
rect 109904 230085 109939 230113
rect 109967 230085 110001 230113
rect 110029 230085 110064 230113
rect 109904 230051 110064 230085
rect 109904 230023 109939 230051
rect 109967 230023 110001 230051
rect 110029 230023 110064 230051
rect 109904 229989 110064 230023
rect 109904 229961 109939 229989
rect 109967 229961 110001 229989
rect 110029 229961 110064 229989
rect 109904 229944 110064 229961
rect 125264 230175 125424 230192
rect 125264 230147 125299 230175
rect 125327 230147 125361 230175
rect 125389 230147 125424 230175
rect 125264 230113 125424 230147
rect 125264 230085 125299 230113
rect 125327 230085 125361 230113
rect 125389 230085 125424 230113
rect 125264 230051 125424 230085
rect 125264 230023 125299 230051
rect 125327 230023 125361 230051
rect 125389 230023 125424 230051
rect 125264 229989 125424 230023
rect 125264 229961 125299 229989
rect 125327 229961 125361 229989
rect 125389 229961 125424 229989
rect 125264 229944 125424 229961
rect 140624 230175 140784 230192
rect 140624 230147 140659 230175
rect 140687 230147 140721 230175
rect 140749 230147 140784 230175
rect 140624 230113 140784 230147
rect 140624 230085 140659 230113
rect 140687 230085 140721 230113
rect 140749 230085 140784 230113
rect 140624 230051 140784 230085
rect 140624 230023 140659 230051
rect 140687 230023 140721 230051
rect 140749 230023 140784 230051
rect 140624 229989 140784 230023
rect 140624 229961 140659 229989
rect 140687 229961 140721 229989
rect 140749 229961 140784 229989
rect 140624 229944 140784 229961
rect 155984 230175 156144 230192
rect 155984 230147 156019 230175
rect 156047 230147 156081 230175
rect 156109 230147 156144 230175
rect 155984 230113 156144 230147
rect 155984 230085 156019 230113
rect 156047 230085 156081 230113
rect 156109 230085 156144 230113
rect 155984 230051 156144 230085
rect 155984 230023 156019 230051
rect 156047 230023 156081 230051
rect 156109 230023 156144 230051
rect 155984 229989 156144 230023
rect 155984 229961 156019 229989
rect 156047 229961 156081 229989
rect 156109 229961 156144 229989
rect 155984 229944 156144 229961
rect 171344 230175 171504 230192
rect 171344 230147 171379 230175
rect 171407 230147 171441 230175
rect 171469 230147 171504 230175
rect 171344 230113 171504 230147
rect 171344 230085 171379 230113
rect 171407 230085 171441 230113
rect 171469 230085 171504 230113
rect 171344 230051 171504 230085
rect 171344 230023 171379 230051
rect 171407 230023 171441 230051
rect 171469 230023 171504 230051
rect 171344 229989 171504 230023
rect 171344 229961 171379 229989
rect 171407 229961 171441 229989
rect 171469 229961 171504 229989
rect 171344 229944 171504 229961
rect 186704 230175 186864 230192
rect 186704 230147 186739 230175
rect 186767 230147 186801 230175
rect 186829 230147 186864 230175
rect 186704 230113 186864 230147
rect 186704 230085 186739 230113
rect 186767 230085 186801 230113
rect 186829 230085 186864 230113
rect 186704 230051 186864 230085
rect 186704 230023 186739 230051
rect 186767 230023 186801 230051
rect 186829 230023 186864 230051
rect 186704 229989 186864 230023
rect 186704 229961 186739 229989
rect 186767 229961 186801 229989
rect 186829 229961 186864 229989
rect 186704 229944 186864 229961
rect 202064 230175 202224 230192
rect 202064 230147 202099 230175
rect 202127 230147 202161 230175
rect 202189 230147 202224 230175
rect 202064 230113 202224 230147
rect 202064 230085 202099 230113
rect 202127 230085 202161 230113
rect 202189 230085 202224 230113
rect 202064 230051 202224 230085
rect 202064 230023 202099 230051
rect 202127 230023 202161 230051
rect 202189 230023 202224 230051
rect 202064 229989 202224 230023
rect 202064 229961 202099 229989
rect 202127 229961 202161 229989
rect 202189 229961 202224 229989
rect 202064 229944 202224 229961
rect 217424 230175 217584 230192
rect 217424 230147 217459 230175
rect 217487 230147 217521 230175
rect 217549 230147 217584 230175
rect 217424 230113 217584 230147
rect 217424 230085 217459 230113
rect 217487 230085 217521 230113
rect 217549 230085 217584 230113
rect 217424 230051 217584 230085
rect 217424 230023 217459 230051
rect 217487 230023 217521 230051
rect 217549 230023 217584 230051
rect 217424 229989 217584 230023
rect 217424 229961 217459 229989
rect 217487 229961 217521 229989
rect 217549 229961 217584 229989
rect 217424 229944 217584 229961
rect 232784 230175 232944 230192
rect 232784 230147 232819 230175
rect 232847 230147 232881 230175
rect 232909 230147 232944 230175
rect 232784 230113 232944 230147
rect 232784 230085 232819 230113
rect 232847 230085 232881 230113
rect 232909 230085 232944 230113
rect 232784 230051 232944 230085
rect 232784 230023 232819 230051
rect 232847 230023 232881 230051
rect 232909 230023 232944 230051
rect 232784 229989 232944 230023
rect 232784 229961 232819 229989
rect 232847 229961 232881 229989
rect 232909 229961 232944 229989
rect 232784 229944 232944 229961
rect 248144 230175 248304 230192
rect 248144 230147 248179 230175
rect 248207 230147 248241 230175
rect 248269 230147 248304 230175
rect 248144 230113 248304 230147
rect 248144 230085 248179 230113
rect 248207 230085 248241 230113
rect 248269 230085 248304 230113
rect 248144 230051 248304 230085
rect 248144 230023 248179 230051
rect 248207 230023 248241 230051
rect 248269 230023 248304 230051
rect 248144 229989 248304 230023
rect 248144 229961 248179 229989
rect 248207 229961 248241 229989
rect 248269 229961 248304 229989
rect 248144 229944 248304 229961
rect 263504 230175 263664 230192
rect 263504 230147 263539 230175
rect 263567 230147 263601 230175
rect 263629 230147 263664 230175
rect 263504 230113 263664 230147
rect 263504 230085 263539 230113
rect 263567 230085 263601 230113
rect 263629 230085 263664 230113
rect 263504 230051 263664 230085
rect 263504 230023 263539 230051
rect 263567 230023 263601 230051
rect 263629 230023 263664 230051
rect 263504 229989 263664 230023
rect 263504 229961 263539 229989
rect 263567 229961 263601 229989
rect 263629 229961 263664 229989
rect 263504 229944 263664 229961
rect 278864 230175 279024 230192
rect 278864 230147 278899 230175
rect 278927 230147 278961 230175
rect 278989 230147 279024 230175
rect 278864 230113 279024 230147
rect 278864 230085 278899 230113
rect 278927 230085 278961 230113
rect 278989 230085 279024 230113
rect 278864 230051 279024 230085
rect 278864 230023 278899 230051
rect 278927 230023 278961 230051
rect 278989 230023 279024 230051
rect 278864 229989 279024 230023
rect 278864 229961 278899 229989
rect 278927 229961 278961 229989
rect 278989 229961 279024 229989
rect 278864 229944 279024 229961
rect 102224 227175 102384 227192
rect 102224 227147 102259 227175
rect 102287 227147 102321 227175
rect 102349 227147 102384 227175
rect 102224 227113 102384 227147
rect 102224 227085 102259 227113
rect 102287 227085 102321 227113
rect 102349 227085 102384 227113
rect 102224 227051 102384 227085
rect 102224 227023 102259 227051
rect 102287 227023 102321 227051
rect 102349 227023 102384 227051
rect 102224 226989 102384 227023
rect 102224 226961 102259 226989
rect 102287 226961 102321 226989
rect 102349 226961 102384 226989
rect 102224 226944 102384 226961
rect 117584 227175 117744 227192
rect 117584 227147 117619 227175
rect 117647 227147 117681 227175
rect 117709 227147 117744 227175
rect 117584 227113 117744 227147
rect 117584 227085 117619 227113
rect 117647 227085 117681 227113
rect 117709 227085 117744 227113
rect 117584 227051 117744 227085
rect 117584 227023 117619 227051
rect 117647 227023 117681 227051
rect 117709 227023 117744 227051
rect 117584 226989 117744 227023
rect 117584 226961 117619 226989
rect 117647 226961 117681 226989
rect 117709 226961 117744 226989
rect 117584 226944 117744 226961
rect 132944 227175 133104 227192
rect 132944 227147 132979 227175
rect 133007 227147 133041 227175
rect 133069 227147 133104 227175
rect 132944 227113 133104 227147
rect 132944 227085 132979 227113
rect 133007 227085 133041 227113
rect 133069 227085 133104 227113
rect 132944 227051 133104 227085
rect 132944 227023 132979 227051
rect 133007 227023 133041 227051
rect 133069 227023 133104 227051
rect 132944 226989 133104 227023
rect 132944 226961 132979 226989
rect 133007 226961 133041 226989
rect 133069 226961 133104 226989
rect 132944 226944 133104 226961
rect 148304 227175 148464 227192
rect 148304 227147 148339 227175
rect 148367 227147 148401 227175
rect 148429 227147 148464 227175
rect 148304 227113 148464 227147
rect 148304 227085 148339 227113
rect 148367 227085 148401 227113
rect 148429 227085 148464 227113
rect 148304 227051 148464 227085
rect 148304 227023 148339 227051
rect 148367 227023 148401 227051
rect 148429 227023 148464 227051
rect 148304 226989 148464 227023
rect 148304 226961 148339 226989
rect 148367 226961 148401 226989
rect 148429 226961 148464 226989
rect 148304 226944 148464 226961
rect 163664 227175 163824 227192
rect 163664 227147 163699 227175
rect 163727 227147 163761 227175
rect 163789 227147 163824 227175
rect 163664 227113 163824 227147
rect 163664 227085 163699 227113
rect 163727 227085 163761 227113
rect 163789 227085 163824 227113
rect 163664 227051 163824 227085
rect 163664 227023 163699 227051
rect 163727 227023 163761 227051
rect 163789 227023 163824 227051
rect 163664 226989 163824 227023
rect 163664 226961 163699 226989
rect 163727 226961 163761 226989
rect 163789 226961 163824 226989
rect 163664 226944 163824 226961
rect 179024 227175 179184 227192
rect 179024 227147 179059 227175
rect 179087 227147 179121 227175
rect 179149 227147 179184 227175
rect 179024 227113 179184 227147
rect 179024 227085 179059 227113
rect 179087 227085 179121 227113
rect 179149 227085 179184 227113
rect 179024 227051 179184 227085
rect 179024 227023 179059 227051
rect 179087 227023 179121 227051
rect 179149 227023 179184 227051
rect 179024 226989 179184 227023
rect 179024 226961 179059 226989
rect 179087 226961 179121 226989
rect 179149 226961 179184 226989
rect 179024 226944 179184 226961
rect 194384 227175 194544 227192
rect 194384 227147 194419 227175
rect 194447 227147 194481 227175
rect 194509 227147 194544 227175
rect 194384 227113 194544 227147
rect 194384 227085 194419 227113
rect 194447 227085 194481 227113
rect 194509 227085 194544 227113
rect 194384 227051 194544 227085
rect 194384 227023 194419 227051
rect 194447 227023 194481 227051
rect 194509 227023 194544 227051
rect 194384 226989 194544 227023
rect 194384 226961 194419 226989
rect 194447 226961 194481 226989
rect 194509 226961 194544 226989
rect 194384 226944 194544 226961
rect 209744 227175 209904 227192
rect 209744 227147 209779 227175
rect 209807 227147 209841 227175
rect 209869 227147 209904 227175
rect 209744 227113 209904 227147
rect 209744 227085 209779 227113
rect 209807 227085 209841 227113
rect 209869 227085 209904 227113
rect 209744 227051 209904 227085
rect 209744 227023 209779 227051
rect 209807 227023 209841 227051
rect 209869 227023 209904 227051
rect 209744 226989 209904 227023
rect 209744 226961 209779 226989
rect 209807 226961 209841 226989
rect 209869 226961 209904 226989
rect 209744 226944 209904 226961
rect 225104 227175 225264 227192
rect 225104 227147 225139 227175
rect 225167 227147 225201 227175
rect 225229 227147 225264 227175
rect 225104 227113 225264 227147
rect 225104 227085 225139 227113
rect 225167 227085 225201 227113
rect 225229 227085 225264 227113
rect 225104 227051 225264 227085
rect 225104 227023 225139 227051
rect 225167 227023 225201 227051
rect 225229 227023 225264 227051
rect 225104 226989 225264 227023
rect 225104 226961 225139 226989
rect 225167 226961 225201 226989
rect 225229 226961 225264 226989
rect 225104 226944 225264 226961
rect 240464 227175 240624 227192
rect 240464 227147 240499 227175
rect 240527 227147 240561 227175
rect 240589 227147 240624 227175
rect 240464 227113 240624 227147
rect 240464 227085 240499 227113
rect 240527 227085 240561 227113
rect 240589 227085 240624 227113
rect 240464 227051 240624 227085
rect 240464 227023 240499 227051
rect 240527 227023 240561 227051
rect 240589 227023 240624 227051
rect 240464 226989 240624 227023
rect 240464 226961 240499 226989
rect 240527 226961 240561 226989
rect 240589 226961 240624 226989
rect 240464 226944 240624 226961
rect 255824 227175 255984 227192
rect 255824 227147 255859 227175
rect 255887 227147 255921 227175
rect 255949 227147 255984 227175
rect 255824 227113 255984 227147
rect 255824 227085 255859 227113
rect 255887 227085 255921 227113
rect 255949 227085 255984 227113
rect 255824 227051 255984 227085
rect 255824 227023 255859 227051
rect 255887 227023 255921 227051
rect 255949 227023 255984 227051
rect 255824 226989 255984 227023
rect 255824 226961 255859 226989
rect 255887 226961 255921 226989
rect 255949 226961 255984 226989
rect 255824 226944 255984 226961
rect 271184 227175 271344 227192
rect 271184 227147 271219 227175
rect 271247 227147 271281 227175
rect 271309 227147 271344 227175
rect 271184 227113 271344 227147
rect 271184 227085 271219 227113
rect 271247 227085 271281 227113
rect 271309 227085 271344 227113
rect 271184 227051 271344 227085
rect 271184 227023 271219 227051
rect 271247 227023 271281 227051
rect 271309 227023 271344 227051
rect 271184 226989 271344 227023
rect 271184 226961 271219 226989
rect 271247 226961 271281 226989
rect 271309 226961 271344 226989
rect 271184 226944 271344 226961
rect 279189 227175 279499 235961
rect 279189 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 279499 227175
rect 279189 227113 279499 227147
rect 279189 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 279499 227113
rect 279189 227051 279499 227085
rect 279189 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 279499 227051
rect 279189 226989 279499 227023
rect 279189 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 279499 226989
rect 109904 221175 110064 221192
rect 109904 221147 109939 221175
rect 109967 221147 110001 221175
rect 110029 221147 110064 221175
rect 109904 221113 110064 221147
rect 109904 221085 109939 221113
rect 109967 221085 110001 221113
rect 110029 221085 110064 221113
rect 109904 221051 110064 221085
rect 109904 221023 109939 221051
rect 109967 221023 110001 221051
rect 110029 221023 110064 221051
rect 109904 220989 110064 221023
rect 109904 220961 109939 220989
rect 109967 220961 110001 220989
rect 110029 220961 110064 220989
rect 109904 220944 110064 220961
rect 125264 221175 125424 221192
rect 125264 221147 125299 221175
rect 125327 221147 125361 221175
rect 125389 221147 125424 221175
rect 125264 221113 125424 221147
rect 125264 221085 125299 221113
rect 125327 221085 125361 221113
rect 125389 221085 125424 221113
rect 125264 221051 125424 221085
rect 125264 221023 125299 221051
rect 125327 221023 125361 221051
rect 125389 221023 125424 221051
rect 125264 220989 125424 221023
rect 125264 220961 125299 220989
rect 125327 220961 125361 220989
rect 125389 220961 125424 220989
rect 125264 220944 125424 220961
rect 140624 221175 140784 221192
rect 140624 221147 140659 221175
rect 140687 221147 140721 221175
rect 140749 221147 140784 221175
rect 140624 221113 140784 221147
rect 140624 221085 140659 221113
rect 140687 221085 140721 221113
rect 140749 221085 140784 221113
rect 140624 221051 140784 221085
rect 140624 221023 140659 221051
rect 140687 221023 140721 221051
rect 140749 221023 140784 221051
rect 140624 220989 140784 221023
rect 140624 220961 140659 220989
rect 140687 220961 140721 220989
rect 140749 220961 140784 220989
rect 140624 220944 140784 220961
rect 155984 221175 156144 221192
rect 155984 221147 156019 221175
rect 156047 221147 156081 221175
rect 156109 221147 156144 221175
rect 155984 221113 156144 221147
rect 155984 221085 156019 221113
rect 156047 221085 156081 221113
rect 156109 221085 156144 221113
rect 155984 221051 156144 221085
rect 155984 221023 156019 221051
rect 156047 221023 156081 221051
rect 156109 221023 156144 221051
rect 155984 220989 156144 221023
rect 155984 220961 156019 220989
rect 156047 220961 156081 220989
rect 156109 220961 156144 220989
rect 155984 220944 156144 220961
rect 171344 221175 171504 221192
rect 171344 221147 171379 221175
rect 171407 221147 171441 221175
rect 171469 221147 171504 221175
rect 171344 221113 171504 221147
rect 171344 221085 171379 221113
rect 171407 221085 171441 221113
rect 171469 221085 171504 221113
rect 171344 221051 171504 221085
rect 171344 221023 171379 221051
rect 171407 221023 171441 221051
rect 171469 221023 171504 221051
rect 171344 220989 171504 221023
rect 171344 220961 171379 220989
rect 171407 220961 171441 220989
rect 171469 220961 171504 220989
rect 171344 220944 171504 220961
rect 186704 221175 186864 221192
rect 186704 221147 186739 221175
rect 186767 221147 186801 221175
rect 186829 221147 186864 221175
rect 186704 221113 186864 221147
rect 186704 221085 186739 221113
rect 186767 221085 186801 221113
rect 186829 221085 186864 221113
rect 186704 221051 186864 221085
rect 186704 221023 186739 221051
rect 186767 221023 186801 221051
rect 186829 221023 186864 221051
rect 186704 220989 186864 221023
rect 186704 220961 186739 220989
rect 186767 220961 186801 220989
rect 186829 220961 186864 220989
rect 186704 220944 186864 220961
rect 202064 221175 202224 221192
rect 202064 221147 202099 221175
rect 202127 221147 202161 221175
rect 202189 221147 202224 221175
rect 202064 221113 202224 221147
rect 202064 221085 202099 221113
rect 202127 221085 202161 221113
rect 202189 221085 202224 221113
rect 202064 221051 202224 221085
rect 202064 221023 202099 221051
rect 202127 221023 202161 221051
rect 202189 221023 202224 221051
rect 202064 220989 202224 221023
rect 202064 220961 202099 220989
rect 202127 220961 202161 220989
rect 202189 220961 202224 220989
rect 202064 220944 202224 220961
rect 217424 221175 217584 221192
rect 217424 221147 217459 221175
rect 217487 221147 217521 221175
rect 217549 221147 217584 221175
rect 217424 221113 217584 221147
rect 217424 221085 217459 221113
rect 217487 221085 217521 221113
rect 217549 221085 217584 221113
rect 217424 221051 217584 221085
rect 217424 221023 217459 221051
rect 217487 221023 217521 221051
rect 217549 221023 217584 221051
rect 217424 220989 217584 221023
rect 217424 220961 217459 220989
rect 217487 220961 217521 220989
rect 217549 220961 217584 220989
rect 217424 220944 217584 220961
rect 232784 221175 232944 221192
rect 232784 221147 232819 221175
rect 232847 221147 232881 221175
rect 232909 221147 232944 221175
rect 232784 221113 232944 221147
rect 232784 221085 232819 221113
rect 232847 221085 232881 221113
rect 232909 221085 232944 221113
rect 232784 221051 232944 221085
rect 232784 221023 232819 221051
rect 232847 221023 232881 221051
rect 232909 221023 232944 221051
rect 232784 220989 232944 221023
rect 232784 220961 232819 220989
rect 232847 220961 232881 220989
rect 232909 220961 232944 220989
rect 232784 220944 232944 220961
rect 248144 221175 248304 221192
rect 248144 221147 248179 221175
rect 248207 221147 248241 221175
rect 248269 221147 248304 221175
rect 248144 221113 248304 221147
rect 248144 221085 248179 221113
rect 248207 221085 248241 221113
rect 248269 221085 248304 221113
rect 248144 221051 248304 221085
rect 248144 221023 248179 221051
rect 248207 221023 248241 221051
rect 248269 221023 248304 221051
rect 248144 220989 248304 221023
rect 248144 220961 248179 220989
rect 248207 220961 248241 220989
rect 248269 220961 248304 220989
rect 248144 220944 248304 220961
rect 263504 221175 263664 221192
rect 263504 221147 263539 221175
rect 263567 221147 263601 221175
rect 263629 221147 263664 221175
rect 263504 221113 263664 221147
rect 263504 221085 263539 221113
rect 263567 221085 263601 221113
rect 263629 221085 263664 221113
rect 263504 221051 263664 221085
rect 263504 221023 263539 221051
rect 263567 221023 263601 221051
rect 263629 221023 263664 221051
rect 263504 220989 263664 221023
rect 263504 220961 263539 220989
rect 263567 220961 263601 220989
rect 263629 220961 263664 220989
rect 263504 220944 263664 220961
rect 278864 221175 279024 221192
rect 278864 221147 278899 221175
rect 278927 221147 278961 221175
rect 278989 221147 279024 221175
rect 278864 221113 279024 221147
rect 278864 221085 278899 221113
rect 278927 221085 278961 221113
rect 278989 221085 279024 221113
rect 278864 221051 279024 221085
rect 278864 221023 278899 221051
rect 278927 221023 278961 221051
rect 278989 221023 279024 221051
rect 278864 220989 279024 221023
rect 278864 220961 278899 220989
rect 278927 220961 278961 220989
rect 278989 220961 279024 220989
rect 278864 220944 279024 220961
rect 102224 218175 102384 218192
rect 102224 218147 102259 218175
rect 102287 218147 102321 218175
rect 102349 218147 102384 218175
rect 102224 218113 102384 218147
rect 102224 218085 102259 218113
rect 102287 218085 102321 218113
rect 102349 218085 102384 218113
rect 102224 218051 102384 218085
rect 102224 218023 102259 218051
rect 102287 218023 102321 218051
rect 102349 218023 102384 218051
rect 102224 217989 102384 218023
rect 102224 217961 102259 217989
rect 102287 217961 102321 217989
rect 102349 217961 102384 217989
rect 102224 217944 102384 217961
rect 117584 218175 117744 218192
rect 117584 218147 117619 218175
rect 117647 218147 117681 218175
rect 117709 218147 117744 218175
rect 117584 218113 117744 218147
rect 117584 218085 117619 218113
rect 117647 218085 117681 218113
rect 117709 218085 117744 218113
rect 117584 218051 117744 218085
rect 117584 218023 117619 218051
rect 117647 218023 117681 218051
rect 117709 218023 117744 218051
rect 117584 217989 117744 218023
rect 117584 217961 117619 217989
rect 117647 217961 117681 217989
rect 117709 217961 117744 217989
rect 117584 217944 117744 217961
rect 132944 218175 133104 218192
rect 132944 218147 132979 218175
rect 133007 218147 133041 218175
rect 133069 218147 133104 218175
rect 132944 218113 133104 218147
rect 132944 218085 132979 218113
rect 133007 218085 133041 218113
rect 133069 218085 133104 218113
rect 132944 218051 133104 218085
rect 132944 218023 132979 218051
rect 133007 218023 133041 218051
rect 133069 218023 133104 218051
rect 132944 217989 133104 218023
rect 132944 217961 132979 217989
rect 133007 217961 133041 217989
rect 133069 217961 133104 217989
rect 132944 217944 133104 217961
rect 148304 218175 148464 218192
rect 148304 218147 148339 218175
rect 148367 218147 148401 218175
rect 148429 218147 148464 218175
rect 148304 218113 148464 218147
rect 148304 218085 148339 218113
rect 148367 218085 148401 218113
rect 148429 218085 148464 218113
rect 148304 218051 148464 218085
rect 148304 218023 148339 218051
rect 148367 218023 148401 218051
rect 148429 218023 148464 218051
rect 148304 217989 148464 218023
rect 148304 217961 148339 217989
rect 148367 217961 148401 217989
rect 148429 217961 148464 217989
rect 148304 217944 148464 217961
rect 163664 218175 163824 218192
rect 163664 218147 163699 218175
rect 163727 218147 163761 218175
rect 163789 218147 163824 218175
rect 163664 218113 163824 218147
rect 163664 218085 163699 218113
rect 163727 218085 163761 218113
rect 163789 218085 163824 218113
rect 163664 218051 163824 218085
rect 163664 218023 163699 218051
rect 163727 218023 163761 218051
rect 163789 218023 163824 218051
rect 163664 217989 163824 218023
rect 163664 217961 163699 217989
rect 163727 217961 163761 217989
rect 163789 217961 163824 217989
rect 163664 217944 163824 217961
rect 179024 218175 179184 218192
rect 179024 218147 179059 218175
rect 179087 218147 179121 218175
rect 179149 218147 179184 218175
rect 179024 218113 179184 218147
rect 179024 218085 179059 218113
rect 179087 218085 179121 218113
rect 179149 218085 179184 218113
rect 179024 218051 179184 218085
rect 179024 218023 179059 218051
rect 179087 218023 179121 218051
rect 179149 218023 179184 218051
rect 179024 217989 179184 218023
rect 179024 217961 179059 217989
rect 179087 217961 179121 217989
rect 179149 217961 179184 217989
rect 179024 217944 179184 217961
rect 194384 218175 194544 218192
rect 194384 218147 194419 218175
rect 194447 218147 194481 218175
rect 194509 218147 194544 218175
rect 194384 218113 194544 218147
rect 194384 218085 194419 218113
rect 194447 218085 194481 218113
rect 194509 218085 194544 218113
rect 194384 218051 194544 218085
rect 194384 218023 194419 218051
rect 194447 218023 194481 218051
rect 194509 218023 194544 218051
rect 194384 217989 194544 218023
rect 194384 217961 194419 217989
rect 194447 217961 194481 217989
rect 194509 217961 194544 217989
rect 194384 217944 194544 217961
rect 209744 218175 209904 218192
rect 209744 218147 209779 218175
rect 209807 218147 209841 218175
rect 209869 218147 209904 218175
rect 209744 218113 209904 218147
rect 209744 218085 209779 218113
rect 209807 218085 209841 218113
rect 209869 218085 209904 218113
rect 209744 218051 209904 218085
rect 209744 218023 209779 218051
rect 209807 218023 209841 218051
rect 209869 218023 209904 218051
rect 209744 217989 209904 218023
rect 209744 217961 209779 217989
rect 209807 217961 209841 217989
rect 209869 217961 209904 217989
rect 209744 217944 209904 217961
rect 225104 218175 225264 218192
rect 225104 218147 225139 218175
rect 225167 218147 225201 218175
rect 225229 218147 225264 218175
rect 225104 218113 225264 218147
rect 225104 218085 225139 218113
rect 225167 218085 225201 218113
rect 225229 218085 225264 218113
rect 225104 218051 225264 218085
rect 225104 218023 225139 218051
rect 225167 218023 225201 218051
rect 225229 218023 225264 218051
rect 225104 217989 225264 218023
rect 225104 217961 225139 217989
rect 225167 217961 225201 217989
rect 225229 217961 225264 217989
rect 225104 217944 225264 217961
rect 240464 218175 240624 218192
rect 240464 218147 240499 218175
rect 240527 218147 240561 218175
rect 240589 218147 240624 218175
rect 240464 218113 240624 218147
rect 240464 218085 240499 218113
rect 240527 218085 240561 218113
rect 240589 218085 240624 218113
rect 240464 218051 240624 218085
rect 240464 218023 240499 218051
rect 240527 218023 240561 218051
rect 240589 218023 240624 218051
rect 240464 217989 240624 218023
rect 240464 217961 240499 217989
rect 240527 217961 240561 217989
rect 240589 217961 240624 217989
rect 240464 217944 240624 217961
rect 255824 218175 255984 218192
rect 255824 218147 255859 218175
rect 255887 218147 255921 218175
rect 255949 218147 255984 218175
rect 255824 218113 255984 218147
rect 255824 218085 255859 218113
rect 255887 218085 255921 218113
rect 255949 218085 255984 218113
rect 255824 218051 255984 218085
rect 255824 218023 255859 218051
rect 255887 218023 255921 218051
rect 255949 218023 255984 218051
rect 255824 217989 255984 218023
rect 255824 217961 255859 217989
rect 255887 217961 255921 217989
rect 255949 217961 255984 217989
rect 255824 217944 255984 217961
rect 271184 218175 271344 218192
rect 271184 218147 271219 218175
rect 271247 218147 271281 218175
rect 271309 218147 271344 218175
rect 271184 218113 271344 218147
rect 271184 218085 271219 218113
rect 271247 218085 271281 218113
rect 271309 218085 271344 218113
rect 271184 218051 271344 218085
rect 271184 218023 271219 218051
rect 271247 218023 271281 218051
rect 271309 218023 271344 218051
rect 271184 217989 271344 218023
rect 271184 217961 271219 217989
rect 271247 217961 271281 217989
rect 271309 217961 271344 217989
rect 271184 217944 271344 217961
rect 279189 218175 279499 226961
rect 279189 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 279499 218175
rect 279189 218113 279499 218147
rect 279189 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 279499 218113
rect 279189 218051 279499 218085
rect 279189 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 279499 218051
rect 279189 217989 279499 218023
rect 279189 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 279499 217989
rect 98966 215866 98994 215871
rect 98854 145385 98882 145390
rect 98910 208474 98938 208479
rect 98798 124217 98826 124222
rect 98854 141946 98882 141951
rect 98742 46601 98770 46606
rect 98798 119770 98826 119775
rect 96729 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 97039 41175
rect 96729 41113 97039 41147
rect 96729 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 97039 41113
rect 96729 41051 97039 41085
rect 96729 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 97039 41051
rect 96729 40989 97039 41023
rect 96729 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 97039 40989
rect 96729 32175 97039 40961
rect 96729 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 97039 32175
rect 96729 32113 97039 32147
rect 96729 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 97039 32113
rect 96729 32051 97039 32085
rect 96729 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 97039 32051
rect 96729 31989 97039 32023
rect 96729 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 97039 31989
rect 96729 23175 97039 31961
rect 96729 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 97039 23175
rect 96729 23113 97039 23147
rect 96729 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 97039 23113
rect 96729 23051 97039 23085
rect 96729 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 97039 23051
rect 96729 22989 97039 23023
rect 96729 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 97039 22989
rect 96729 14175 97039 22961
rect 98798 18410 98826 119742
rect 98854 39578 98882 141918
rect 98910 103082 98938 208446
rect 98966 110138 98994 215838
rect 109904 212175 110064 212192
rect 109904 212147 109939 212175
rect 109967 212147 110001 212175
rect 110029 212147 110064 212175
rect 109904 212113 110064 212147
rect 109904 212085 109939 212113
rect 109967 212085 110001 212113
rect 110029 212085 110064 212113
rect 109904 212051 110064 212085
rect 109904 212023 109939 212051
rect 109967 212023 110001 212051
rect 110029 212023 110064 212051
rect 109904 211989 110064 212023
rect 109904 211961 109939 211989
rect 109967 211961 110001 211989
rect 110029 211961 110064 211989
rect 109904 211944 110064 211961
rect 125264 212175 125424 212192
rect 125264 212147 125299 212175
rect 125327 212147 125361 212175
rect 125389 212147 125424 212175
rect 125264 212113 125424 212147
rect 125264 212085 125299 212113
rect 125327 212085 125361 212113
rect 125389 212085 125424 212113
rect 125264 212051 125424 212085
rect 125264 212023 125299 212051
rect 125327 212023 125361 212051
rect 125389 212023 125424 212051
rect 125264 211989 125424 212023
rect 125264 211961 125299 211989
rect 125327 211961 125361 211989
rect 125389 211961 125424 211989
rect 125264 211944 125424 211961
rect 140624 212175 140784 212192
rect 140624 212147 140659 212175
rect 140687 212147 140721 212175
rect 140749 212147 140784 212175
rect 140624 212113 140784 212147
rect 140624 212085 140659 212113
rect 140687 212085 140721 212113
rect 140749 212085 140784 212113
rect 140624 212051 140784 212085
rect 140624 212023 140659 212051
rect 140687 212023 140721 212051
rect 140749 212023 140784 212051
rect 140624 211989 140784 212023
rect 140624 211961 140659 211989
rect 140687 211961 140721 211989
rect 140749 211961 140784 211989
rect 140624 211944 140784 211961
rect 155984 212175 156144 212192
rect 155984 212147 156019 212175
rect 156047 212147 156081 212175
rect 156109 212147 156144 212175
rect 155984 212113 156144 212147
rect 155984 212085 156019 212113
rect 156047 212085 156081 212113
rect 156109 212085 156144 212113
rect 155984 212051 156144 212085
rect 155984 212023 156019 212051
rect 156047 212023 156081 212051
rect 156109 212023 156144 212051
rect 155984 211989 156144 212023
rect 155984 211961 156019 211989
rect 156047 211961 156081 211989
rect 156109 211961 156144 211989
rect 155984 211944 156144 211961
rect 171344 212175 171504 212192
rect 171344 212147 171379 212175
rect 171407 212147 171441 212175
rect 171469 212147 171504 212175
rect 171344 212113 171504 212147
rect 171344 212085 171379 212113
rect 171407 212085 171441 212113
rect 171469 212085 171504 212113
rect 171344 212051 171504 212085
rect 171344 212023 171379 212051
rect 171407 212023 171441 212051
rect 171469 212023 171504 212051
rect 171344 211989 171504 212023
rect 171344 211961 171379 211989
rect 171407 211961 171441 211989
rect 171469 211961 171504 211989
rect 171344 211944 171504 211961
rect 186704 212175 186864 212192
rect 186704 212147 186739 212175
rect 186767 212147 186801 212175
rect 186829 212147 186864 212175
rect 186704 212113 186864 212147
rect 186704 212085 186739 212113
rect 186767 212085 186801 212113
rect 186829 212085 186864 212113
rect 186704 212051 186864 212085
rect 186704 212023 186739 212051
rect 186767 212023 186801 212051
rect 186829 212023 186864 212051
rect 186704 211989 186864 212023
rect 186704 211961 186739 211989
rect 186767 211961 186801 211989
rect 186829 211961 186864 211989
rect 186704 211944 186864 211961
rect 202064 212175 202224 212192
rect 202064 212147 202099 212175
rect 202127 212147 202161 212175
rect 202189 212147 202224 212175
rect 202064 212113 202224 212147
rect 202064 212085 202099 212113
rect 202127 212085 202161 212113
rect 202189 212085 202224 212113
rect 202064 212051 202224 212085
rect 202064 212023 202099 212051
rect 202127 212023 202161 212051
rect 202189 212023 202224 212051
rect 202064 211989 202224 212023
rect 202064 211961 202099 211989
rect 202127 211961 202161 211989
rect 202189 211961 202224 211989
rect 202064 211944 202224 211961
rect 217424 212175 217584 212192
rect 217424 212147 217459 212175
rect 217487 212147 217521 212175
rect 217549 212147 217584 212175
rect 217424 212113 217584 212147
rect 217424 212085 217459 212113
rect 217487 212085 217521 212113
rect 217549 212085 217584 212113
rect 217424 212051 217584 212085
rect 217424 212023 217459 212051
rect 217487 212023 217521 212051
rect 217549 212023 217584 212051
rect 217424 211989 217584 212023
rect 217424 211961 217459 211989
rect 217487 211961 217521 211989
rect 217549 211961 217584 211989
rect 217424 211944 217584 211961
rect 232784 212175 232944 212192
rect 232784 212147 232819 212175
rect 232847 212147 232881 212175
rect 232909 212147 232944 212175
rect 232784 212113 232944 212147
rect 232784 212085 232819 212113
rect 232847 212085 232881 212113
rect 232909 212085 232944 212113
rect 232784 212051 232944 212085
rect 232784 212023 232819 212051
rect 232847 212023 232881 212051
rect 232909 212023 232944 212051
rect 232784 211989 232944 212023
rect 232784 211961 232819 211989
rect 232847 211961 232881 211989
rect 232909 211961 232944 211989
rect 232784 211944 232944 211961
rect 248144 212175 248304 212192
rect 248144 212147 248179 212175
rect 248207 212147 248241 212175
rect 248269 212147 248304 212175
rect 248144 212113 248304 212147
rect 248144 212085 248179 212113
rect 248207 212085 248241 212113
rect 248269 212085 248304 212113
rect 248144 212051 248304 212085
rect 248144 212023 248179 212051
rect 248207 212023 248241 212051
rect 248269 212023 248304 212051
rect 248144 211989 248304 212023
rect 248144 211961 248179 211989
rect 248207 211961 248241 211989
rect 248269 211961 248304 211989
rect 248144 211944 248304 211961
rect 263504 212175 263664 212192
rect 263504 212147 263539 212175
rect 263567 212147 263601 212175
rect 263629 212147 263664 212175
rect 263504 212113 263664 212147
rect 263504 212085 263539 212113
rect 263567 212085 263601 212113
rect 263629 212085 263664 212113
rect 263504 212051 263664 212085
rect 263504 212023 263539 212051
rect 263567 212023 263601 212051
rect 263629 212023 263664 212051
rect 263504 211989 263664 212023
rect 263504 211961 263539 211989
rect 263567 211961 263601 211989
rect 263629 211961 263664 211989
rect 263504 211944 263664 211961
rect 278864 212175 279024 212192
rect 278864 212147 278899 212175
rect 278927 212147 278961 212175
rect 278989 212147 279024 212175
rect 278864 212113 279024 212147
rect 278864 212085 278899 212113
rect 278927 212085 278961 212113
rect 278989 212085 279024 212113
rect 278864 212051 279024 212085
rect 278864 212023 278899 212051
rect 278927 212023 278961 212051
rect 278989 212023 279024 212051
rect 278864 211989 279024 212023
rect 278864 211961 278899 211989
rect 278927 211961 278961 211989
rect 278989 211961 279024 211989
rect 278864 211944 279024 211961
rect 102224 209175 102384 209192
rect 102224 209147 102259 209175
rect 102287 209147 102321 209175
rect 102349 209147 102384 209175
rect 102224 209113 102384 209147
rect 102224 209085 102259 209113
rect 102287 209085 102321 209113
rect 102349 209085 102384 209113
rect 102224 209051 102384 209085
rect 102224 209023 102259 209051
rect 102287 209023 102321 209051
rect 102349 209023 102384 209051
rect 102224 208989 102384 209023
rect 102224 208961 102259 208989
rect 102287 208961 102321 208989
rect 102349 208961 102384 208989
rect 102224 208944 102384 208961
rect 117584 209175 117744 209192
rect 117584 209147 117619 209175
rect 117647 209147 117681 209175
rect 117709 209147 117744 209175
rect 117584 209113 117744 209147
rect 117584 209085 117619 209113
rect 117647 209085 117681 209113
rect 117709 209085 117744 209113
rect 117584 209051 117744 209085
rect 117584 209023 117619 209051
rect 117647 209023 117681 209051
rect 117709 209023 117744 209051
rect 117584 208989 117744 209023
rect 117584 208961 117619 208989
rect 117647 208961 117681 208989
rect 117709 208961 117744 208989
rect 117584 208944 117744 208961
rect 132944 209175 133104 209192
rect 132944 209147 132979 209175
rect 133007 209147 133041 209175
rect 133069 209147 133104 209175
rect 132944 209113 133104 209147
rect 132944 209085 132979 209113
rect 133007 209085 133041 209113
rect 133069 209085 133104 209113
rect 132944 209051 133104 209085
rect 132944 209023 132979 209051
rect 133007 209023 133041 209051
rect 133069 209023 133104 209051
rect 132944 208989 133104 209023
rect 132944 208961 132979 208989
rect 133007 208961 133041 208989
rect 133069 208961 133104 208989
rect 132944 208944 133104 208961
rect 148304 209175 148464 209192
rect 148304 209147 148339 209175
rect 148367 209147 148401 209175
rect 148429 209147 148464 209175
rect 148304 209113 148464 209147
rect 148304 209085 148339 209113
rect 148367 209085 148401 209113
rect 148429 209085 148464 209113
rect 148304 209051 148464 209085
rect 148304 209023 148339 209051
rect 148367 209023 148401 209051
rect 148429 209023 148464 209051
rect 148304 208989 148464 209023
rect 148304 208961 148339 208989
rect 148367 208961 148401 208989
rect 148429 208961 148464 208989
rect 148304 208944 148464 208961
rect 163664 209175 163824 209192
rect 163664 209147 163699 209175
rect 163727 209147 163761 209175
rect 163789 209147 163824 209175
rect 163664 209113 163824 209147
rect 163664 209085 163699 209113
rect 163727 209085 163761 209113
rect 163789 209085 163824 209113
rect 163664 209051 163824 209085
rect 163664 209023 163699 209051
rect 163727 209023 163761 209051
rect 163789 209023 163824 209051
rect 163664 208989 163824 209023
rect 163664 208961 163699 208989
rect 163727 208961 163761 208989
rect 163789 208961 163824 208989
rect 163664 208944 163824 208961
rect 179024 209175 179184 209192
rect 179024 209147 179059 209175
rect 179087 209147 179121 209175
rect 179149 209147 179184 209175
rect 179024 209113 179184 209147
rect 179024 209085 179059 209113
rect 179087 209085 179121 209113
rect 179149 209085 179184 209113
rect 179024 209051 179184 209085
rect 179024 209023 179059 209051
rect 179087 209023 179121 209051
rect 179149 209023 179184 209051
rect 179024 208989 179184 209023
rect 179024 208961 179059 208989
rect 179087 208961 179121 208989
rect 179149 208961 179184 208989
rect 179024 208944 179184 208961
rect 194384 209175 194544 209192
rect 194384 209147 194419 209175
rect 194447 209147 194481 209175
rect 194509 209147 194544 209175
rect 194384 209113 194544 209147
rect 194384 209085 194419 209113
rect 194447 209085 194481 209113
rect 194509 209085 194544 209113
rect 194384 209051 194544 209085
rect 194384 209023 194419 209051
rect 194447 209023 194481 209051
rect 194509 209023 194544 209051
rect 194384 208989 194544 209023
rect 194384 208961 194419 208989
rect 194447 208961 194481 208989
rect 194509 208961 194544 208989
rect 194384 208944 194544 208961
rect 209744 209175 209904 209192
rect 209744 209147 209779 209175
rect 209807 209147 209841 209175
rect 209869 209147 209904 209175
rect 209744 209113 209904 209147
rect 209744 209085 209779 209113
rect 209807 209085 209841 209113
rect 209869 209085 209904 209113
rect 209744 209051 209904 209085
rect 209744 209023 209779 209051
rect 209807 209023 209841 209051
rect 209869 209023 209904 209051
rect 209744 208989 209904 209023
rect 209744 208961 209779 208989
rect 209807 208961 209841 208989
rect 209869 208961 209904 208989
rect 209744 208944 209904 208961
rect 225104 209175 225264 209192
rect 225104 209147 225139 209175
rect 225167 209147 225201 209175
rect 225229 209147 225264 209175
rect 225104 209113 225264 209147
rect 225104 209085 225139 209113
rect 225167 209085 225201 209113
rect 225229 209085 225264 209113
rect 225104 209051 225264 209085
rect 225104 209023 225139 209051
rect 225167 209023 225201 209051
rect 225229 209023 225264 209051
rect 225104 208989 225264 209023
rect 225104 208961 225139 208989
rect 225167 208961 225201 208989
rect 225229 208961 225264 208989
rect 225104 208944 225264 208961
rect 240464 209175 240624 209192
rect 240464 209147 240499 209175
rect 240527 209147 240561 209175
rect 240589 209147 240624 209175
rect 240464 209113 240624 209147
rect 240464 209085 240499 209113
rect 240527 209085 240561 209113
rect 240589 209085 240624 209113
rect 240464 209051 240624 209085
rect 240464 209023 240499 209051
rect 240527 209023 240561 209051
rect 240589 209023 240624 209051
rect 240464 208989 240624 209023
rect 240464 208961 240499 208989
rect 240527 208961 240561 208989
rect 240589 208961 240624 208989
rect 240464 208944 240624 208961
rect 255824 209175 255984 209192
rect 255824 209147 255859 209175
rect 255887 209147 255921 209175
rect 255949 209147 255984 209175
rect 255824 209113 255984 209147
rect 255824 209085 255859 209113
rect 255887 209085 255921 209113
rect 255949 209085 255984 209113
rect 255824 209051 255984 209085
rect 255824 209023 255859 209051
rect 255887 209023 255921 209051
rect 255949 209023 255984 209051
rect 255824 208989 255984 209023
rect 255824 208961 255859 208989
rect 255887 208961 255921 208989
rect 255949 208961 255984 208989
rect 255824 208944 255984 208961
rect 271184 209175 271344 209192
rect 271184 209147 271219 209175
rect 271247 209147 271281 209175
rect 271309 209147 271344 209175
rect 271184 209113 271344 209147
rect 271184 209085 271219 209113
rect 271247 209085 271281 209113
rect 271309 209085 271344 209113
rect 271184 209051 271344 209085
rect 271184 209023 271219 209051
rect 271247 209023 271281 209051
rect 271309 209023 271344 209051
rect 271184 208989 271344 209023
rect 271184 208961 271219 208989
rect 271247 208961 271281 208989
rect 271309 208961 271344 208989
rect 271184 208944 271344 208961
rect 279189 209175 279499 217961
rect 279189 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 279499 209175
rect 279189 209113 279499 209147
rect 279189 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 279499 209113
rect 279189 209051 279499 209085
rect 279189 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 279499 209051
rect 279189 208989 279499 209023
rect 279189 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 279499 208989
rect 109904 203175 110064 203192
rect 109904 203147 109939 203175
rect 109967 203147 110001 203175
rect 110029 203147 110064 203175
rect 109904 203113 110064 203147
rect 109904 203085 109939 203113
rect 109967 203085 110001 203113
rect 110029 203085 110064 203113
rect 109904 203051 110064 203085
rect 109904 203023 109939 203051
rect 109967 203023 110001 203051
rect 110029 203023 110064 203051
rect 109904 202989 110064 203023
rect 109904 202961 109939 202989
rect 109967 202961 110001 202989
rect 110029 202961 110064 202989
rect 109904 202944 110064 202961
rect 125264 203175 125424 203192
rect 125264 203147 125299 203175
rect 125327 203147 125361 203175
rect 125389 203147 125424 203175
rect 125264 203113 125424 203147
rect 125264 203085 125299 203113
rect 125327 203085 125361 203113
rect 125389 203085 125424 203113
rect 125264 203051 125424 203085
rect 125264 203023 125299 203051
rect 125327 203023 125361 203051
rect 125389 203023 125424 203051
rect 125264 202989 125424 203023
rect 125264 202961 125299 202989
rect 125327 202961 125361 202989
rect 125389 202961 125424 202989
rect 125264 202944 125424 202961
rect 140624 203175 140784 203192
rect 140624 203147 140659 203175
rect 140687 203147 140721 203175
rect 140749 203147 140784 203175
rect 140624 203113 140784 203147
rect 140624 203085 140659 203113
rect 140687 203085 140721 203113
rect 140749 203085 140784 203113
rect 140624 203051 140784 203085
rect 140624 203023 140659 203051
rect 140687 203023 140721 203051
rect 140749 203023 140784 203051
rect 140624 202989 140784 203023
rect 140624 202961 140659 202989
rect 140687 202961 140721 202989
rect 140749 202961 140784 202989
rect 140624 202944 140784 202961
rect 155984 203175 156144 203192
rect 155984 203147 156019 203175
rect 156047 203147 156081 203175
rect 156109 203147 156144 203175
rect 155984 203113 156144 203147
rect 155984 203085 156019 203113
rect 156047 203085 156081 203113
rect 156109 203085 156144 203113
rect 155984 203051 156144 203085
rect 155984 203023 156019 203051
rect 156047 203023 156081 203051
rect 156109 203023 156144 203051
rect 155984 202989 156144 203023
rect 155984 202961 156019 202989
rect 156047 202961 156081 202989
rect 156109 202961 156144 202989
rect 155984 202944 156144 202961
rect 171344 203175 171504 203192
rect 171344 203147 171379 203175
rect 171407 203147 171441 203175
rect 171469 203147 171504 203175
rect 171344 203113 171504 203147
rect 171344 203085 171379 203113
rect 171407 203085 171441 203113
rect 171469 203085 171504 203113
rect 171344 203051 171504 203085
rect 171344 203023 171379 203051
rect 171407 203023 171441 203051
rect 171469 203023 171504 203051
rect 171344 202989 171504 203023
rect 171344 202961 171379 202989
rect 171407 202961 171441 202989
rect 171469 202961 171504 202989
rect 171344 202944 171504 202961
rect 186704 203175 186864 203192
rect 186704 203147 186739 203175
rect 186767 203147 186801 203175
rect 186829 203147 186864 203175
rect 186704 203113 186864 203147
rect 186704 203085 186739 203113
rect 186767 203085 186801 203113
rect 186829 203085 186864 203113
rect 186704 203051 186864 203085
rect 186704 203023 186739 203051
rect 186767 203023 186801 203051
rect 186829 203023 186864 203051
rect 186704 202989 186864 203023
rect 186704 202961 186739 202989
rect 186767 202961 186801 202989
rect 186829 202961 186864 202989
rect 186704 202944 186864 202961
rect 202064 203175 202224 203192
rect 202064 203147 202099 203175
rect 202127 203147 202161 203175
rect 202189 203147 202224 203175
rect 202064 203113 202224 203147
rect 202064 203085 202099 203113
rect 202127 203085 202161 203113
rect 202189 203085 202224 203113
rect 202064 203051 202224 203085
rect 202064 203023 202099 203051
rect 202127 203023 202161 203051
rect 202189 203023 202224 203051
rect 202064 202989 202224 203023
rect 202064 202961 202099 202989
rect 202127 202961 202161 202989
rect 202189 202961 202224 202989
rect 202064 202944 202224 202961
rect 217424 203175 217584 203192
rect 217424 203147 217459 203175
rect 217487 203147 217521 203175
rect 217549 203147 217584 203175
rect 217424 203113 217584 203147
rect 217424 203085 217459 203113
rect 217487 203085 217521 203113
rect 217549 203085 217584 203113
rect 217424 203051 217584 203085
rect 217424 203023 217459 203051
rect 217487 203023 217521 203051
rect 217549 203023 217584 203051
rect 217424 202989 217584 203023
rect 217424 202961 217459 202989
rect 217487 202961 217521 202989
rect 217549 202961 217584 202989
rect 217424 202944 217584 202961
rect 232784 203175 232944 203192
rect 232784 203147 232819 203175
rect 232847 203147 232881 203175
rect 232909 203147 232944 203175
rect 232784 203113 232944 203147
rect 232784 203085 232819 203113
rect 232847 203085 232881 203113
rect 232909 203085 232944 203113
rect 232784 203051 232944 203085
rect 232784 203023 232819 203051
rect 232847 203023 232881 203051
rect 232909 203023 232944 203051
rect 232784 202989 232944 203023
rect 232784 202961 232819 202989
rect 232847 202961 232881 202989
rect 232909 202961 232944 202989
rect 232784 202944 232944 202961
rect 248144 203175 248304 203192
rect 248144 203147 248179 203175
rect 248207 203147 248241 203175
rect 248269 203147 248304 203175
rect 248144 203113 248304 203147
rect 248144 203085 248179 203113
rect 248207 203085 248241 203113
rect 248269 203085 248304 203113
rect 248144 203051 248304 203085
rect 248144 203023 248179 203051
rect 248207 203023 248241 203051
rect 248269 203023 248304 203051
rect 248144 202989 248304 203023
rect 248144 202961 248179 202989
rect 248207 202961 248241 202989
rect 248269 202961 248304 202989
rect 248144 202944 248304 202961
rect 263504 203175 263664 203192
rect 263504 203147 263539 203175
rect 263567 203147 263601 203175
rect 263629 203147 263664 203175
rect 263504 203113 263664 203147
rect 263504 203085 263539 203113
rect 263567 203085 263601 203113
rect 263629 203085 263664 203113
rect 263504 203051 263664 203085
rect 263504 203023 263539 203051
rect 263567 203023 263601 203051
rect 263629 203023 263664 203051
rect 263504 202989 263664 203023
rect 263504 202961 263539 202989
rect 263567 202961 263601 202989
rect 263629 202961 263664 202989
rect 263504 202944 263664 202961
rect 278864 203175 279024 203192
rect 278864 203147 278899 203175
rect 278927 203147 278961 203175
rect 278989 203147 279024 203175
rect 278864 203113 279024 203147
rect 278864 203085 278899 203113
rect 278927 203085 278961 203113
rect 278989 203085 279024 203113
rect 278864 203051 279024 203085
rect 278864 203023 278899 203051
rect 278927 203023 278961 203051
rect 278989 203023 279024 203051
rect 278864 202989 279024 203023
rect 278864 202961 278899 202989
rect 278927 202961 278961 202989
rect 278989 202961 279024 202989
rect 278864 202944 279024 202961
rect 102224 200175 102384 200192
rect 102224 200147 102259 200175
rect 102287 200147 102321 200175
rect 102349 200147 102384 200175
rect 102224 200113 102384 200147
rect 102224 200085 102259 200113
rect 102287 200085 102321 200113
rect 102349 200085 102384 200113
rect 102224 200051 102384 200085
rect 102224 200023 102259 200051
rect 102287 200023 102321 200051
rect 102349 200023 102384 200051
rect 102224 199989 102384 200023
rect 102224 199961 102259 199989
rect 102287 199961 102321 199989
rect 102349 199961 102384 199989
rect 102224 199944 102384 199961
rect 117584 200175 117744 200192
rect 117584 200147 117619 200175
rect 117647 200147 117681 200175
rect 117709 200147 117744 200175
rect 117584 200113 117744 200147
rect 117584 200085 117619 200113
rect 117647 200085 117681 200113
rect 117709 200085 117744 200113
rect 117584 200051 117744 200085
rect 117584 200023 117619 200051
rect 117647 200023 117681 200051
rect 117709 200023 117744 200051
rect 117584 199989 117744 200023
rect 117584 199961 117619 199989
rect 117647 199961 117681 199989
rect 117709 199961 117744 199989
rect 117584 199944 117744 199961
rect 132944 200175 133104 200192
rect 132944 200147 132979 200175
rect 133007 200147 133041 200175
rect 133069 200147 133104 200175
rect 132944 200113 133104 200147
rect 132944 200085 132979 200113
rect 133007 200085 133041 200113
rect 133069 200085 133104 200113
rect 132944 200051 133104 200085
rect 132944 200023 132979 200051
rect 133007 200023 133041 200051
rect 133069 200023 133104 200051
rect 132944 199989 133104 200023
rect 132944 199961 132979 199989
rect 133007 199961 133041 199989
rect 133069 199961 133104 199989
rect 132944 199944 133104 199961
rect 148304 200175 148464 200192
rect 148304 200147 148339 200175
rect 148367 200147 148401 200175
rect 148429 200147 148464 200175
rect 148304 200113 148464 200147
rect 148304 200085 148339 200113
rect 148367 200085 148401 200113
rect 148429 200085 148464 200113
rect 148304 200051 148464 200085
rect 148304 200023 148339 200051
rect 148367 200023 148401 200051
rect 148429 200023 148464 200051
rect 148304 199989 148464 200023
rect 148304 199961 148339 199989
rect 148367 199961 148401 199989
rect 148429 199961 148464 199989
rect 148304 199944 148464 199961
rect 163664 200175 163824 200192
rect 163664 200147 163699 200175
rect 163727 200147 163761 200175
rect 163789 200147 163824 200175
rect 163664 200113 163824 200147
rect 163664 200085 163699 200113
rect 163727 200085 163761 200113
rect 163789 200085 163824 200113
rect 163664 200051 163824 200085
rect 163664 200023 163699 200051
rect 163727 200023 163761 200051
rect 163789 200023 163824 200051
rect 163664 199989 163824 200023
rect 163664 199961 163699 199989
rect 163727 199961 163761 199989
rect 163789 199961 163824 199989
rect 163664 199944 163824 199961
rect 179024 200175 179184 200192
rect 179024 200147 179059 200175
rect 179087 200147 179121 200175
rect 179149 200147 179184 200175
rect 179024 200113 179184 200147
rect 179024 200085 179059 200113
rect 179087 200085 179121 200113
rect 179149 200085 179184 200113
rect 179024 200051 179184 200085
rect 179024 200023 179059 200051
rect 179087 200023 179121 200051
rect 179149 200023 179184 200051
rect 179024 199989 179184 200023
rect 179024 199961 179059 199989
rect 179087 199961 179121 199989
rect 179149 199961 179184 199989
rect 179024 199944 179184 199961
rect 194384 200175 194544 200192
rect 194384 200147 194419 200175
rect 194447 200147 194481 200175
rect 194509 200147 194544 200175
rect 194384 200113 194544 200147
rect 194384 200085 194419 200113
rect 194447 200085 194481 200113
rect 194509 200085 194544 200113
rect 194384 200051 194544 200085
rect 194384 200023 194419 200051
rect 194447 200023 194481 200051
rect 194509 200023 194544 200051
rect 194384 199989 194544 200023
rect 194384 199961 194419 199989
rect 194447 199961 194481 199989
rect 194509 199961 194544 199989
rect 194384 199944 194544 199961
rect 209744 200175 209904 200192
rect 209744 200147 209779 200175
rect 209807 200147 209841 200175
rect 209869 200147 209904 200175
rect 209744 200113 209904 200147
rect 209744 200085 209779 200113
rect 209807 200085 209841 200113
rect 209869 200085 209904 200113
rect 209744 200051 209904 200085
rect 209744 200023 209779 200051
rect 209807 200023 209841 200051
rect 209869 200023 209904 200051
rect 209744 199989 209904 200023
rect 209744 199961 209779 199989
rect 209807 199961 209841 199989
rect 209869 199961 209904 199989
rect 209744 199944 209904 199961
rect 225104 200175 225264 200192
rect 225104 200147 225139 200175
rect 225167 200147 225201 200175
rect 225229 200147 225264 200175
rect 225104 200113 225264 200147
rect 225104 200085 225139 200113
rect 225167 200085 225201 200113
rect 225229 200085 225264 200113
rect 225104 200051 225264 200085
rect 225104 200023 225139 200051
rect 225167 200023 225201 200051
rect 225229 200023 225264 200051
rect 225104 199989 225264 200023
rect 225104 199961 225139 199989
rect 225167 199961 225201 199989
rect 225229 199961 225264 199989
rect 225104 199944 225264 199961
rect 240464 200175 240624 200192
rect 240464 200147 240499 200175
rect 240527 200147 240561 200175
rect 240589 200147 240624 200175
rect 240464 200113 240624 200147
rect 240464 200085 240499 200113
rect 240527 200085 240561 200113
rect 240589 200085 240624 200113
rect 240464 200051 240624 200085
rect 240464 200023 240499 200051
rect 240527 200023 240561 200051
rect 240589 200023 240624 200051
rect 240464 199989 240624 200023
rect 240464 199961 240499 199989
rect 240527 199961 240561 199989
rect 240589 199961 240624 199989
rect 240464 199944 240624 199961
rect 255824 200175 255984 200192
rect 255824 200147 255859 200175
rect 255887 200147 255921 200175
rect 255949 200147 255984 200175
rect 255824 200113 255984 200147
rect 255824 200085 255859 200113
rect 255887 200085 255921 200113
rect 255949 200085 255984 200113
rect 255824 200051 255984 200085
rect 255824 200023 255859 200051
rect 255887 200023 255921 200051
rect 255949 200023 255984 200051
rect 255824 199989 255984 200023
rect 255824 199961 255859 199989
rect 255887 199961 255921 199989
rect 255949 199961 255984 199989
rect 255824 199944 255984 199961
rect 271184 200175 271344 200192
rect 271184 200147 271219 200175
rect 271247 200147 271281 200175
rect 271309 200147 271344 200175
rect 271184 200113 271344 200147
rect 271184 200085 271219 200113
rect 271247 200085 271281 200113
rect 271309 200085 271344 200113
rect 271184 200051 271344 200085
rect 271184 200023 271219 200051
rect 271247 200023 271281 200051
rect 271309 200023 271344 200051
rect 271184 199989 271344 200023
rect 271184 199961 271219 199989
rect 271247 199961 271281 199989
rect 271309 199961 271344 199989
rect 271184 199944 271344 199961
rect 279189 200175 279499 208961
rect 279189 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 279499 200175
rect 279189 200113 279499 200147
rect 279189 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 279499 200113
rect 279189 200051 279499 200085
rect 279189 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 279499 200051
rect 279189 199989 279499 200023
rect 279189 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 279499 199989
rect 109904 194175 110064 194192
rect 109904 194147 109939 194175
rect 109967 194147 110001 194175
rect 110029 194147 110064 194175
rect 109904 194113 110064 194147
rect 109904 194085 109939 194113
rect 109967 194085 110001 194113
rect 110029 194085 110064 194113
rect 109904 194051 110064 194085
rect 109904 194023 109939 194051
rect 109967 194023 110001 194051
rect 110029 194023 110064 194051
rect 109904 193989 110064 194023
rect 109904 193961 109939 193989
rect 109967 193961 110001 193989
rect 110029 193961 110064 193989
rect 109904 193944 110064 193961
rect 125264 194175 125424 194192
rect 125264 194147 125299 194175
rect 125327 194147 125361 194175
rect 125389 194147 125424 194175
rect 125264 194113 125424 194147
rect 125264 194085 125299 194113
rect 125327 194085 125361 194113
rect 125389 194085 125424 194113
rect 125264 194051 125424 194085
rect 125264 194023 125299 194051
rect 125327 194023 125361 194051
rect 125389 194023 125424 194051
rect 125264 193989 125424 194023
rect 125264 193961 125299 193989
rect 125327 193961 125361 193989
rect 125389 193961 125424 193989
rect 125264 193944 125424 193961
rect 140624 194175 140784 194192
rect 140624 194147 140659 194175
rect 140687 194147 140721 194175
rect 140749 194147 140784 194175
rect 140624 194113 140784 194147
rect 140624 194085 140659 194113
rect 140687 194085 140721 194113
rect 140749 194085 140784 194113
rect 140624 194051 140784 194085
rect 140624 194023 140659 194051
rect 140687 194023 140721 194051
rect 140749 194023 140784 194051
rect 140624 193989 140784 194023
rect 140624 193961 140659 193989
rect 140687 193961 140721 193989
rect 140749 193961 140784 193989
rect 140624 193944 140784 193961
rect 155984 194175 156144 194192
rect 155984 194147 156019 194175
rect 156047 194147 156081 194175
rect 156109 194147 156144 194175
rect 155984 194113 156144 194147
rect 155984 194085 156019 194113
rect 156047 194085 156081 194113
rect 156109 194085 156144 194113
rect 155984 194051 156144 194085
rect 155984 194023 156019 194051
rect 156047 194023 156081 194051
rect 156109 194023 156144 194051
rect 155984 193989 156144 194023
rect 155984 193961 156019 193989
rect 156047 193961 156081 193989
rect 156109 193961 156144 193989
rect 155984 193944 156144 193961
rect 171344 194175 171504 194192
rect 171344 194147 171379 194175
rect 171407 194147 171441 194175
rect 171469 194147 171504 194175
rect 171344 194113 171504 194147
rect 171344 194085 171379 194113
rect 171407 194085 171441 194113
rect 171469 194085 171504 194113
rect 171344 194051 171504 194085
rect 171344 194023 171379 194051
rect 171407 194023 171441 194051
rect 171469 194023 171504 194051
rect 171344 193989 171504 194023
rect 171344 193961 171379 193989
rect 171407 193961 171441 193989
rect 171469 193961 171504 193989
rect 171344 193944 171504 193961
rect 186704 194175 186864 194192
rect 186704 194147 186739 194175
rect 186767 194147 186801 194175
rect 186829 194147 186864 194175
rect 186704 194113 186864 194147
rect 186704 194085 186739 194113
rect 186767 194085 186801 194113
rect 186829 194085 186864 194113
rect 186704 194051 186864 194085
rect 186704 194023 186739 194051
rect 186767 194023 186801 194051
rect 186829 194023 186864 194051
rect 186704 193989 186864 194023
rect 186704 193961 186739 193989
rect 186767 193961 186801 193989
rect 186829 193961 186864 193989
rect 186704 193944 186864 193961
rect 202064 194175 202224 194192
rect 202064 194147 202099 194175
rect 202127 194147 202161 194175
rect 202189 194147 202224 194175
rect 202064 194113 202224 194147
rect 202064 194085 202099 194113
rect 202127 194085 202161 194113
rect 202189 194085 202224 194113
rect 202064 194051 202224 194085
rect 202064 194023 202099 194051
rect 202127 194023 202161 194051
rect 202189 194023 202224 194051
rect 202064 193989 202224 194023
rect 202064 193961 202099 193989
rect 202127 193961 202161 193989
rect 202189 193961 202224 193989
rect 202064 193944 202224 193961
rect 217424 194175 217584 194192
rect 217424 194147 217459 194175
rect 217487 194147 217521 194175
rect 217549 194147 217584 194175
rect 217424 194113 217584 194147
rect 217424 194085 217459 194113
rect 217487 194085 217521 194113
rect 217549 194085 217584 194113
rect 217424 194051 217584 194085
rect 217424 194023 217459 194051
rect 217487 194023 217521 194051
rect 217549 194023 217584 194051
rect 217424 193989 217584 194023
rect 217424 193961 217459 193989
rect 217487 193961 217521 193989
rect 217549 193961 217584 193989
rect 217424 193944 217584 193961
rect 232784 194175 232944 194192
rect 232784 194147 232819 194175
rect 232847 194147 232881 194175
rect 232909 194147 232944 194175
rect 232784 194113 232944 194147
rect 232784 194085 232819 194113
rect 232847 194085 232881 194113
rect 232909 194085 232944 194113
rect 232784 194051 232944 194085
rect 232784 194023 232819 194051
rect 232847 194023 232881 194051
rect 232909 194023 232944 194051
rect 232784 193989 232944 194023
rect 232784 193961 232819 193989
rect 232847 193961 232881 193989
rect 232909 193961 232944 193989
rect 232784 193944 232944 193961
rect 248144 194175 248304 194192
rect 248144 194147 248179 194175
rect 248207 194147 248241 194175
rect 248269 194147 248304 194175
rect 248144 194113 248304 194147
rect 248144 194085 248179 194113
rect 248207 194085 248241 194113
rect 248269 194085 248304 194113
rect 248144 194051 248304 194085
rect 248144 194023 248179 194051
rect 248207 194023 248241 194051
rect 248269 194023 248304 194051
rect 248144 193989 248304 194023
rect 248144 193961 248179 193989
rect 248207 193961 248241 193989
rect 248269 193961 248304 193989
rect 248144 193944 248304 193961
rect 263504 194175 263664 194192
rect 263504 194147 263539 194175
rect 263567 194147 263601 194175
rect 263629 194147 263664 194175
rect 263504 194113 263664 194147
rect 263504 194085 263539 194113
rect 263567 194085 263601 194113
rect 263629 194085 263664 194113
rect 263504 194051 263664 194085
rect 263504 194023 263539 194051
rect 263567 194023 263601 194051
rect 263629 194023 263664 194051
rect 263504 193989 263664 194023
rect 263504 193961 263539 193989
rect 263567 193961 263601 193989
rect 263629 193961 263664 193989
rect 263504 193944 263664 193961
rect 278864 194175 279024 194192
rect 278864 194147 278899 194175
rect 278927 194147 278961 194175
rect 278989 194147 279024 194175
rect 278864 194113 279024 194147
rect 278864 194085 278899 194113
rect 278927 194085 278961 194113
rect 278989 194085 279024 194113
rect 278864 194051 279024 194085
rect 278864 194023 278899 194051
rect 278927 194023 278961 194051
rect 278989 194023 279024 194051
rect 278864 193989 279024 194023
rect 278864 193961 278899 193989
rect 278927 193961 278961 193989
rect 278989 193961 279024 193989
rect 278864 193944 279024 193961
rect 98966 110105 98994 110110
rect 99022 193690 99050 193695
rect 98910 103049 98938 103054
rect 99022 88970 99050 193662
rect 102224 191175 102384 191192
rect 102224 191147 102259 191175
rect 102287 191147 102321 191175
rect 102349 191147 102384 191175
rect 102224 191113 102384 191147
rect 102224 191085 102259 191113
rect 102287 191085 102321 191113
rect 102349 191085 102384 191113
rect 102224 191051 102384 191085
rect 102224 191023 102259 191051
rect 102287 191023 102321 191051
rect 102349 191023 102384 191051
rect 102224 190989 102384 191023
rect 102224 190961 102259 190989
rect 102287 190961 102321 190989
rect 102349 190961 102384 190989
rect 102224 190944 102384 190961
rect 117584 191175 117744 191192
rect 117584 191147 117619 191175
rect 117647 191147 117681 191175
rect 117709 191147 117744 191175
rect 117584 191113 117744 191147
rect 117584 191085 117619 191113
rect 117647 191085 117681 191113
rect 117709 191085 117744 191113
rect 117584 191051 117744 191085
rect 117584 191023 117619 191051
rect 117647 191023 117681 191051
rect 117709 191023 117744 191051
rect 117584 190989 117744 191023
rect 117584 190961 117619 190989
rect 117647 190961 117681 190989
rect 117709 190961 117744 190989
rect 117584 190944 117744 190961
rect 132944 191175 133104 191192
rect 132944 191147 132979 191175
rect 133007 191147 133041 191175
rect 133069 191147 133104 191175
rect 132944 191113 133104 191147
rect 132944 191085 132979 191113
rect 133007 191085 133041 191113
rect 133069 191085 133104 191113
rect 132944 191051 133104 191085
rect 132944 191023 132979 191051
rect 133007 191023 133041 191051
rect 133069 191023 133104 191051
rect 132944 190989 133104 191023
rect 132944 190961 132979 190989
rect 133007 190961 133041 190989
rect 133069 190961 133104 190989
rect 132944 190944 133104 190961
rect 148304 191175 148464 191192
rect 148304 191147 148339 191175
rect 148367 191147 148401 191175
rect 148429 191147 148464 191175
rect 148304 191113 148464 191147
rect 148304 191085 148339 191113
rect 148367 191085 148401 191113
rect 148429 191085 148464 191113
rect 148304 191051 148464 191085
rect 148304 191023 148339 191051
rect 148367 191023 148401 191051
rect 148429 191023 148464 191051
rect 148304 190989 148464 191023
rect 148304 190961 148339 190989
rect 148367 190961 148401 190989
rect 148429 190961 148464 190989
rect 148304 190944 148464 190961
rect 163664 191175 163824 191192
rect 163664 191147 163699 191175
rect 163727 191147 163761 191175
rect 163789 191147 163824 191175
rect 163664 191113 163824 191147
rect 163664 191085 163699 191113
rect 163727 191085 163761 191113
rect 163789 191085 163824 191113
rect 163664 191051 163824 191085
rect 163664 191023 163699 191051
rect 163727 191023 163761 191051
rect 163789 191023 163824 191051
rect 163664 190989 163824 191023
rect 163664 190961 163699 190989
rect 163727 190961 163761 190989
rect 163789 190961 163824 190989
rect 163664 190944 163824 190961
rect 179024 191175 179184 191192
rect 179024 191147 179059 191175
rect 179087 191147 179121 191175
rect 179149 191147 179184 191175
rect 179024 191113 179184 191147
rect 179024 191085 179059 191113
rect 179087 191085 179121 191113
rect 179149 191085 179184 191113
rect 179024 191051 179184 191085
rect 179024 191023 179059 191051
rect 179087 191023 179121 191051
rect 179149 191023 179184 191051
rect 179024 190989 179184 191023
rect 179024 190961 179059 190989
rect 179087 190961 179121 190989
rect 179149 190961 179184 190989
rect 179024 190944 179184 190961
rect 194384 191175 194544 191192
rect 194384 191147 194419 191175
rect 194447 191147 194481 191175
rect 194509 191147 194544 191175
rect 194384 191113 194544 191147
rect 194384 191085 194419 191113
rect 194447 191085 194481 191113
rect 194509 191085 194544 191113
rect 194384 191051 194544 191085
rect 194384 191023 194419 191051
rect 194447 191023 194481 191051
rect 194509 191023 194544 191051
rect 194384 190989 194544 191023
rect 194384 190961 194419 190989
rect 194447 190961 194481 190989
rect 194509 190961 194544 190989
rect 194384 190944 194544 190961
rect 209744 191175 209904 191192
rect 209744 191147 209779 191175
rect 209807 191147 209841 191175
rect 209869 191147 209904 191175
rect 209744 191113 209904 191147
rect 209744 191085 209779 191113
rect 209807 191085 209841 191113
rect 209869 191085 209904 191113
rect 209744 191051 209904 191085
rect 209744 191023 209779 191051
rect 209807 191023 209841 191051
rect 209869 191023 209904 191051
rect 209744 190989 209904 191023
rect 209744 190961 209779 190989
rect 209807 190961 209841 190989
rect 209869 190961 209904 190989
rect 209744 190944 209904 190961
rect 225104 191175 225264 191192
rect 225104 191147 225139 191175
rect 225167 191147 225201 191175
rect 225229 191147 225264 191175
rect 225104 191113 225264 191147
rect 225104 191085 225139 191113
rect 225167 191085 225201 191113
rect 225229 191085 225264 191113
rect 225104 191051 225264 191085
rect 225104 191023 225139 191051
rect 225167 191023 225201 191051
rect 225229 191023 225264 191051
rect 225104 190989 225264 191023
rect 225104 190961 225139 190989
rect 225167 190961 225201 190989
rect 225229 190961 225264 190989
rect 225104 190944 225264 190961
rect 240464 191175 240624 191192
rect 240464 191147 240499 191175
rect 240527 191147 240561 191175
rect 240589 191147 240624 191175
rect 240464 191113 240624 191147
rect 240464 191085 240499 191113
rect 240527 191085 240561 191113
rect 240589 191085 240624 191113
rect 240464 191051 240624 191085
rect 240464 191023 240499 191051
rect 240527 191023 240561 191051
rect 240589 191023 240624 191051
rect 240464 190989 240624 191023
rect 240464 190961 240499 190989
rect 240527 190961 240561 190989
rect 240589 190961 240624 190989
rect 240464 190944 240624 190961
rect 255824 191175 255984 191192
rect 255824 191147 255859 191175
rect 255887 191147 255921 191175
rect 255949 191147 255984 191175
rect 255824 191113 255984 191147
rect 255824 191085 255859 191113
rect 255887 191085 255921 191113
rect 255949 191085 255984 191113
rect 255824 191051 255984 191085
rect 255824 191023 255859 191051
rect 255887 191023 255921 191051
rect 255949 191023 255984 191051
rect 255824 190989 255984 191023
rect 255824 190961 255859 190989
rect 255887 190961 255921 190989
rect 255949 190961 255984 190989
rect 255824 190944 255984 190961
rect 271184 191175 271344 191192
rect 271184 191147 271219 191175
rect 271247 191147 271281 191175
rect 271309 191147 271344 191175
rect 271184 191113 271344 191147
rect 271184 191085 271219 191113
rect 271247 191085 271281 191113
rect 271309 191085 271344 191113
rect 271184 191051 271344 191085
rect 271184 191023 271219 191051
rect 271247 191023 271281 191051
rect 271309 191023 271344 191051
rect 271184 190989 271344 191023
rect 271184 190961 271219 190989
rect 271247 190961 271281 190989
rect 271309 190961 271344 190989
rect 271184 190944 271344 190961
rect 279189 191175 279499 199961
rect 279189 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 279499 191175
rect 279189 191113 279499 191147
rect 279189 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 279499 191113
rect 279189 191051 279499 191085
rect 279189 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 279499 191051
rect 279189 190989 279499 191023
rect 279189 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 279499 190989
rect 109904 185175 110064 185192
rect 109904 185147 109939 185175
rect 109967 185147 110001 185175
rect 110029 185147 110064 185175
rect 109904 185113 110064 185147
rect 109904 185085 109939 185113
rect 109967 185085 110001 185113
rect 110029 185085 110064 185113
rect 109904 185051 110064 185085
rect 109904 185023 109939 185051
rect 109967 185023 110001 185051
rect 110029 185023 110064 185051
rect 109904 184989 110064 185023
rect 109904 184961 109939 184989
rect 109967 184961 110001 184989
rect 110029 184961 110064 184989
rect 109904 184944 110064 184961
rect 125264 185175 125424 185192
rect 125264 185147 125299 185175
rect 125327 185147 125361 185175
rect 125389 185147 125424 185175
rect 125264 185113 125424 185147
rect 125264 185085 125299 185113
rect 125327 185085 125361 185113
rect 125389 185085 125424 185113
rect 125264 185051 125424 185085
rect 125264 185023 125299 185051
rect 125327 185023 125361 185051
rect 125389 185023 125424 185051
rect 125264 184989 125424 185023
rect 125264 184961 125299 184989
rect 125327 184961 125361 184989
rect 125389 184961 125424 184989
rect 125264 184944 125424 184961
rect 140624 185175 140784 185192
rect 140624 185147 140659 185175
rect 140687 185147 140721 185175
rect 140749 185147 140784 185175
rect 140624 185113 140784 185147
rect 140624 185085 140659 185113
rect 140687 185085 140721 185113
rect 140749 185085 140784 185113
rect 140624 185051 140784 185085
rect 140624 185023 140659 185051
rect 140687 185023 140721 185051
rect 140749 185023 140784 185051
rect 140624 184989 140784 185023
rect 140624 184961 140659 184989
rect 140687 184961 140721 184989
rect 140749 184961 140784 184989
rect 140624 184944 140784 184961
rect 155984 185175 156144 185192
rect 155984 185147 156019 185175
rect 156047 185147 156081 185175
rect 156109 185147 156144 185175
rect 155984 185113 156144 185147
rect 155984 185085 156019 185113
rect 156047 185085 156081 185113
rect 156109 185085 156144 185113
rect 155984 185051 156144 185085
rect 155984 185023 156019 185051
rect 156047 185023 156081 185051
rect 156109 185023 156144 185051
rect 155984 184989 156144 185023
rect 155984 184961 156019 184989
rect 156047 184961 156081 184989
rect 156109 184961 156144 184989
rect 155984 184944 156144 184961
rect 171344 185175 171504 185192
rect 171344 185147 171379 185175
rect 171407 185147 171441 185175
rect 171469 185147 171504 185175
rect 171344 185113 171504 185147
rect 171344 185085 171379 185113
rect 171407 185085 171441 185113
rect 171469 185085 171504 185113
rect 171344 185051 171504 185085
rect 171344 185023 171379 185051
rect 171407 185023 171441 185051
rect 171469 185023 171504 185051
rect 171344 184989 171504 185023
rect 171344 184961 171379 184989
rect 171407 184961 171441 184989
rect 171469 184961 171504 184989
rect 171344 184944 171504 184961
rect 186704 185175 186864 185192
rect 186704 185147 186739 185175
rect 186767 185147 186801 185175
rect 186829 185147 186864 185175
rect 186704 185113 186864 185147
rect 186704 185085 186739 185113
rect 186767 185085 186801 185113
rect 186829 185085 186864 185113
rect 186704 185051 186864 185085
rect 186704 185023 186739 185051
rect 186767 185023 186801 185051
rect 186829 185023 186864 185051
rect 186704 184989 186864 185023
rect 186704 184961 186739 184989
rect 186767 184961 186801 184989
rect 186829 184961 186864 184989
rect 186704 184944 186864 184961
rect 202064 185175 202224 185192
rect 202064 185147 202099 185175
rect 202127 185147 202161 185175
rect 202189 185147 202224 185175
rect 202064 185113 202224 185147
rect 202064 185085 202099 185113
rect 202127 185085 202161 185113
rect 202189 185085 202224 185113
rect 202064 185051 202224 185085
rect 202064 185023 202099 185051
rect 202127 185023 202161 185051
rect 202189 185023 202224 185051
rect 202064 184989 202224 185023
rect 202064 184961 202099 184989
rect 202127 184961 202161 184989
rect 202189 184961 202224 184989
rect 202064 184944 202224 184961
rect 217424 185175 217584 185192
rect 217424 185147 217459 185175
rect 217487 185147 217521 185175
rect 217549 185147 217584 185175
rect 217424 185113 217584 185147
rect 217424 185085 217459 185113
rect 217487 185085 217521 185113
rect 217549 185085 217584 185113
rect 217424 185051 217584 185085
rect 217424 185023 217459 185051
rect 217487 185023 217521 185051
rect 217549 185023 217584 185051
rect 217424 184989 217584 185023
rect 217424 184961 217459 184989
rect 217487 184961 217521 184989
rect 217549 184961 217584 184989
rect 217424 184944 217584 184961
rect 232784 185175 232944 185192
rect 232784 185147 232819 185175
rect 232847 185147 232881 185175
rect 232909 185147 232944 185175
rect 232784 185113 232944 185147
rect 232784 185085 232819 185113
rect 232847 185085 232881 185113
rect 232909 185085 232944 185113
rect 232784 185051 232944 185085
rect 232784 185023 232819 185051
rect 232847 185023 232881 185051
rect 232909 185023 232944 185051
rect 232784 184989 232944 185023
rect 232784 184961 232819 184989
rect 232847 184961 232881 184989
rect 232909 184961 232944 184989
rect 232784 184944 232944 184961
rect 248144 185175 248304 185192
rect 248144 185147 248179 185175
rect 248207 185147 248241 185175
rect 248269 185147 248304 185175
rect 248144 185113 248304 185147
rect 248144 185085 248179 185113
rect 248207 185085 248241 185113
rect 248269 185085 248304 185113
rect 248144 185051 248304 185085
rect 248144 185023 248179 185051
rect 248207 185023 248241 185051
rect 248269 185023 248304 185051
rect 248144 184989 248304 185023
rect 248144 184961 248179 184989
rect 248207 184961 248241 184989
rect 248269 184961 248304 184989
rect 248144 184944 248304 184961
rect 263504 185175 263664 185192
rect 263504 185147 263539 185175
rect 263567 185147 263601 185175
rect 263629 185147 263664 185175
rect 263504 185113 263664 185147
rect 263504 185085 263539 185113
rect 263567 185085 263601 185113
rect 263629 185085 263664 185113
rect 263504 185051 263664 185085
rect 263504 185023 263539 185051
rect 263567 185023 263601 185051
rect 263629 185023 263664 185051
rect 263504 184989 263664 185023
rect 263504 184961 263539 184989
rect 263567 184961 263601 184989
rect 263629 184961 263664 184989
rect 263504 184944 263664 184961
rect 278864 185175 279024 185192
rect 278864 185147 278899 185175
rect 278927 185147 278961 185175
rect 278989 185147 279024 185175
rect 278864 185113 279024 185147
rect 278864 185085 278899 185113
rect 278927 185085 278961 185113
rect 278989 185085 279024 185113
rect 278864 185051 279024 185085
rect 278864 185023 278899 185051
rect 278927 185023 278961 185051
rect 278989 185023 279024 185051
rect 278864 184989 279024 185023
rect 278864 184961 278899 184989
rect 278927 184961 278961 184989
rect 278989 184961 279024 184989
rect 278864 184944 279024 184961
rect 102224 182175 102384 182192
rect 102224 182147 102259 182175
rect 102287 182147 102321 182175
rect 102349 182147 102384 182175
rect 102224 182113 102384 182147
rect 102224 182085 102259 182113
rect 102287 182085 102321 182113
rect 102349 182085 102384 182113
rect 102224 182051 102384 182085
rect 102224 182023 102259 182051
rect 102287 182023 102321 182051
rect 102349 182023 102384 182051
rect 102224 181989 102384 182023
rect 102224 181961 102259 181989
rect 102287 181961 102321 181989
rect 102349 181961 102384 181989
rect 102224 181944 102384 181961
rect 117584 182175 117744 182192
rect 117584 182147 117619 182175
rect 117647 182147 117681 182175
rect 117709 182147 117744 182175
rect 117584 182113 117744 182147
rect 117584 182085 117619 182113
rect 117647 182085 117681 182113
rect 117709 182085 117744 182113
rect 117584 182051 117744 182085
rect 117584 182023 117619 182051
rect 117647 182023 117681 182051
rect 117709 182023 117744 182051
rect 117584 181989 117744 182023
rect 117584 181961 117619 181989
rect 117647 181961 117681 181989
rect 117709 181961 117744 181989
rect 117584 181944 117744 181961
rect 132944 182175 133104 182192
rect 132944 182147 132979 182175
rect 133007 182147 133041 182175
rect 133069 182147 133104 182175
rect 132944 182113 133104 182147
rect 132944 182085 132979 182113
rect 133007 182085 133041 182113
rect 133069 182085 133104 182113
rect 132944 182051 133104 182085
rect 132944 182023 132979 182051
rect 133007 182023 133041 182051
rect 133069 182023 133104 182051
rect 132944 181989 133104 182023
rect 132944 181961 132979 181989
rect 133007 181961 133041 181989
rect 133069 181961 133104 181989
rect 132944 181944 133104 181961
rect 148304 182175 148464 182192
rect 148304 182147 148339 182175
rect 148367 182147 148401 182175
rect 148429 182147 148464 182175
rect 148304 182113 148464 182147
rect 148304 182085 148339 182113
rect 148367 182085 148401 182113
rect 148429 182085 148464 182113
rect 148304 182051 148464 182085
rect 148304 182023 148339 182051
rect 148367 182023 148401 182051
rect 148429 182023 148464 182051
rect 148304 181989 148464 182023
rect 148304 181961 148339 181989
rect 148367 181961 148401 181989
rect 148429 181961 148464 181989
rect 148304 181944 148464 181961
rect 163664 182175 163824 182192
rect 163664 182147 163699 182175
rect 163727 182147 163761 182175
rect 163789 182147 163824 182175
rect 163664 182113 163824 182147
rect 163664 182085 163699 182113
rect 163727 182085 163761 182113
rect 163789 182085 163824 182113
rect 163664 182051 163824 182085
rect 163664 182023 163699 182051
rect 163727 182023 163761 182051
rect 163789 182023 163824 182051
rect 163664 181989 163824 182023
rect 163664 181961 163699 181989
rect 163727 181961 163761 181989
rect 163789 181961 163824 181989
rect 163664 181944 163824 181961
rect 179024 182175 179184 182192
rect 179024 182147 179059 182175
rect 179087 182147 179121 182175
rect 179149 182147 179184 182175
rect 179024 182113 179184 182147
rect 179024 182085 179059 182113
rect 179087 182085 179121 182113
rect 179149 182085 179184 182113
rect 179024 182051 179184 182085
rect 179024 182023 179059 182051
rect 179087 182023 179121 182051
rect 179149 182023 179184 182051
rect 179024 181989 179184 182023
rect 179024 181961 179059 181989
rect 179087 181961 179121 181989
rect 179149 181961 179184 181989
rect 179024 181944 179184 181961
rect 194384 182175 194544 182192
rect 194384 182147 194419 182175
rect 194447 182147 194481 182175
rect 194509 182147 194544 182175
rect 194384 182113 194544 182147
rect 194384 182085 194419 182113
rect 194447 182085 194481 182113
rect 194509 182085 194544 182113
rect 194384 182051 194544 182085
rect 194384 182023 194419 182051
rect 194447 182023 194481 182051
rect 194509 182023 194544 182051
rect 194384 181989 194544 182023
rect 194384 181961 194419 181989
rect 194447 181961 194481 181989
rect 194509 181961 194544 181989
rect 194384 181944 194544 181961
rect 209744 182175 209904 182192
rect 209744 182147 209779 182175
rect 209807 182147 209841 182175
rect 209869 182147 209904 182175
rect 209744 182113 209904 182147
rect 209744 182085 209779 182113
rect 209807 182085 209841 182113
rect 209869 182085 209904 182113
rect 209744 182051 209904 182085
rect 209744 182023 209779 182051
rect 209807 182023 209841 182051
rect 209869 182023 209904 182051
rect 209744 181989 209904 182023
rect 209744 181961 209779 181989
rect 209807 181961 209841 181989
rect 209869 181961 209904 181989
rect 209744 181944 209904 181961
rect 225104 182175 225264 182192
rect 225104 182147 225139 182175
rect 225167 182147 225201 182175
rect 225229 182147 225264 182175
rect 225104 182113 225264 182147
rect 225104 182085 225139 182113
rect 225167 182085 225201 182113
rect 225229 182085 225264 182113
rect 225104 182051 225264 182085
rect 225104 182023 225139 182051
rect 225167 182023 225201 182051
rect 225229 182023 225264 182051
rect 225104 181989 225264 182023
rect 225104 181961 225139 181989
rect 225167 181961 225201 181989
rect 225229 181961 225264 181989
rect 225104 181944 225264 181961
rect 240464 182175 240624 182192
rect 240464 182147 240499 182175
rect 240527 182147 240561 182175
rect 240589 182147 240624 182175
rect 240464 182113 240624 182147
rect 240464 182085 240499 182113
rect 240527 182085 240561 182113
rect 240589 182085 240624 182113
rect 240464 182051 240624 182085
rect 240464 182023 240499 182051
rect 240527 182023 240561 182051
rect 240589 182023 240624 182051
rect 240464 181989 240624 182023
rect 240464 181961 240499 181989
rect 240527 181961 240561 181989
rect 240589 181961 240624 181989
rect 240464 181944 240624 181961
rect 255824 182175 255984 182192
rect 255824 182147 255859 182175
rect 255887 182147 255921 182175
rect 255949 182147 255984 182175
rect 255824 182113 255984 182147
rect 255824 182085 255859 182113
rect 255887 182085 255921 182113
rect 255949 182085 255984 182113
rect 255824 182051 255984 182085
rect 255824 182023 255859 182051
rect 255887 182023 255921 182051
rect 255949 182023 255984 182051
rect 255824 181989 255984 182023
rect 255824 181961 255859 181989
rect 255887 181961 255921 181989
rect 255949 181961 255984 181989
rect 255824 181944 255984 181961
rect 271184 182175 271344 182192
rect 271184 182147 271219 182175
rect 271247 182147 271281 182175
rect 271309 182147 271344 182175
rect 271184 182113 271344 182147
rect 271184 182085 271219 182113
rect 271247 182085 271281 182113
rect 271309 182085 271344 182113
rect 271184 182051 271344 182085
rect 271184 182023 271219 182051
rect 271247 182023 271281 182051
rect 271309 182023 271344 182051
rect 271184 181989 271344 182023
rect 271184 181961 271219 181989
rect 271247 181961 271281 181989
rect 271309 181961 271344 181989
rect 271184 181944 271344 181961
rect 279189 182175 279499 190961
rect 279189 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 279499 182175
rect 279189 182113 279499 182147
rect 279189 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 279499 182113
rect 279189 182051 279499 182085
rect 279189 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 279499 182051
rect 279189 181989 279499 182023
rect 279189 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 279499 181989
rect 109904 176175 110064 176192
rect 109904 176147 109939 176175
rect 109967 176147 110001 176175
rect 110029 176147 110064 176175
rect 109904 176113 110064 176147
rect 109904 176085 109939 176113
rect 109967 176085 110001 176113
rect 110029 176085 110064 176113
rect 109904 176051 110064 176085
rect 109904 176023 109939 176051
rect 109967 176023 110001 176051
rect 110029 176023 110064 176051
rect 109904 175989 110064 176023
rect 109904 175961 109939 175989
rect 109967 175961 110001 175989
rect 110029 175961 110064 175989
rect 109904 175944 110064 175961
rect 125264 176175 125424 176192
rect 125264 176147 125299 176175
rect 125327 176147 125361 176175
rect 125389 176147 125424 176175
rect 125264 176113 125424 176147
rect 125264 176085 125299 176113
rect 125327 176085 125361 176113
rect 125389 176085 125424 176113
rect 125264 176051 125424 176085
rect 125264 176023 125299 176051
rect 125327 176023 125361 176051
rect 125389 176023 125424 176051
rect 125264 175989 125424 176023
rect 125264 175961 125299 175989
rect 125327 175961 125361 175989
rect 125389 175961 125424 175989
rect 125264 175944 125424 175961
rect 140624 176175 140784 176192
rect 140624 176147 140659 176175
rect 140687 176147 140721 176175
rect 140749 176147 140784 176175
rect 140624 176113 140784 176147
rect 140624 176085 140659 176113
rect 140687 176085 140721 176113
rect 140749 176085 140784 176113
rect 140624 176051 140784 176085
rect 140624 176023 140659 176051
rect 140687 176023 140721 176051
rect 140749 176023 140784 176051
rect 140624 175989 140784 176023
rect 140624 175961 140659 175989
rect 140687 175961 140721 175989
rect 140749 175961 140784 175989
rect 140624 175944 140784 175961
rect 155984 176175 156144 176192
rect 155984 176147 156019 176175
rect 156047 176147 156081 176175
rect 156109 176147 156144 176175
rect 155984 176113 156144 176147
rect 155984 176085 156019 176113
rect 156047 176085 156081 176113
rect 156109 176085 156144 176113
rect 155984 176051 156144 176085
rect 155984 176023 156019 176051
rect 156047 176023 156081 176051
rect 156109 176023 156144 176051
rect 155984 175989 156144 176023
rect 155984 175961 156019 175989
rect 156047 175961 156081 175989
rect 156109 175961 156144 175989
rect 155984 175944 156144 175961
rect 171344 176175 171504 176192
rect 171344 176147 171379 176175
rect 171407 176147 171441 176175
rect 171469 176147 171504 176175
rect 171344 176113 171504 176147
rect 171344 176085 171379 176113
rect 171407 176085 171441 176113
rect 171469 176085 171504 176113
rect 171344 176051 171504 176085
rect 171344 176023 171379 176051
rect 171407 176023 171441 176051
rect 171469 176023 171504 176051
rect 171344 175989 171504 176023
rect 171344 175961 171379 175989
rect 171407 175961 171441 175989
rect 171469 175961 171504 175989
rect 171344 175944 171504 175961
rect 186704 176175 186864 176192
rect 186704 176147 186739 176175
rect 186767 176147 186801 176175
rect 186829 176147 186864 176175
rect 186704 176113 186864 176147
rect 186704 176085 186739 176113
rect 186767 176085 186801 176113
rect 186829 176085 186864 176113
rect 186704 176051 186864 176085
rect 186704 176023 186739 176051
rect 186767 176023 186801 176051
rect 186829 176023 186864 176051
rect 186704 175989 186864 176023
rect 186704 175961 186739 175989
rect 186767 175961 186801 175989
rect 186829 175961 186864 175989
rect 186704 175944 186864 175961
rect 202064 176175 202224 176192
rect 202064 176147 202099 176175
rect 202127 176147 202161 176175
rect 202189 176147 202224 176175
rect 202064 176113 202224 176147
rect 202064 176085 202099 176113
rect 202127 176085 202161 176113
rect 202189 176085 202224 176113
rect 202064 176051 202224 176085
rect 202064 176023 202099 176051
rect 202127 176023 202161 176051
rect 202189 176023 202224 176051
rect 202064 175989 202224 176023
rect 202064 175961 202099 175989
rect 202127 175961 202161 175989
rect 202189 175961 202224 175989
rect 202064 175944 202224 175961
rect 217424 176175 217584 176192
rect 217424 176147 217459 176175
rect 217487 176147 217521 176175
rect 217549 176147 217584 176175
rect 217424 176113 217584 176147
rect 217424 176085 217459 176113
rect 217487 176085 217521 176113
rect 217549 176085 217584 176113
rect 217424 176051 217584 176085
rect 217424 176023 217459 176051
rect 217487 176023 217521 176051
rect 217549 176023 217584 176051
rect 217424 175989 217584 176023
rect 217424 175961 217459 175989
rect 217487 175961 217521 175989
rect 217549 175961 217584 175989
rect 217424 175944 217584 175961
rect 232784 176175 232944 176192
rect 232784 176147 232819 176175
rect 232847 176147 232881 176175
rect 232909 176147 232944 176175
rect 232784 176113 232944 176147
rect 232784 176085 232819 176113
rect 232847 176085 232881 176113
rect 232909 176085 232944 176113
rect 232784 176051 232944 176085
rect 232784 176023 232819 176051
rect 232847 176023 232881 176051
rect 232909 176023 232944 176051
rect 232784 175989 232944 176023
rect 232784 175961 232819 175989
rect 232847 175961 232881 175989
rect 232909 175961 232944 175989
rect 232784 175944 232944 175961
rect 248144 176175 248304 176192
rect 248144 176147 248179 176175
rect 248207 176147 248241 176175
rect 248269 176147 248304 176175
rect 248144 176113 248304 176147
rect 248144 176085 248179 176113
rect 248207 176085 248241 176113
rect 248269 176085 248304 176113
rect 248144 176051 248304 176085
rect 248144 176023 248179 176051
rect 248207 176023 248241 176051
rect 248269 176023 248304 176051
rect 248144 175989 248304 176023
rect 248144 175961 248179 175989
rect 248207 175961 248241 175989
rect 248269 175961 248304 175989
rect 248144 175944 248304 175961
rect 263504 176175 263664 176192
rect 263504 176147 263539 176175
rect 263567 176147 263601 176175
rect 263629 176147 263664 176175
rect 263504 176113 263664 176147
rect 263504 176085 263539 176113
rect 263567 176085 263601 176113
rect 263629 176085 263664 176113
rect 263504 176051 263664 176085
rect 263504 176023 263539 176051
rect 263567 176023 263601 176051
rect 263629 176023 263664 176051
rect 263504 175989 263664 176023
rect 263504 175961 263539 175989
rect 263567 175961 263601 175989
rect 263629 175961 263664 175989
rect 263504 175944 263664 175961
rect 278864 176175 279024 176192
rect 278864 176147 278899 176175
rect 278927 176147 278961 176175
rect 278989 176147 279024 176175
rect 278864 176113 279024 176147
rect 278864 176085 278899 176113
rect 278927 176085 278961 176113
rect 278989 176085 279024 176113
rect 278864 176051 279024 176085
rect 278864 176023 278899 176051
rect 278927 176023 278961 176051
rect 278989 176023 279024 176051
rect 278864 175989 279024 176023
rect 278864 175961 278899 175989
rect 278927 175961 278961 175989
rect 278989 175961 279024 175989
rect 278864 175944 279024 175961
rect 102224 173175 102384 173192
rect 102224 173147 102259 173175
rect 102287 173147 102321 173175
rect 102349 173147 102384 173175
rect 102224 173113 102384 173147
rect 102224 173085 102259 173113
rect 102287 173085 102321 173113
rect 102349 173085 102384 173113
rect 102224 173051 102384 173085
rect 102224 173023 102259 173051
rect 102287 173023 102321 173051
rect 102349 173023 102384 173051
rect 102224 172989 102384 173023
rect 102224 172961 102259 172989
rect 102287 172961 102321 172989
rect 102349 172961 102384 172989
rect 102224 172944 102384 172961
rect 117584 173175 117744 173192
rect 117584 173147 117619 173175
rect 117647 173147 117681 173175
rect 117709 173147 117744 173175
rect 117584 173113 117744 173147
rect 117584 173085 117619 173113
rect 117647 173085 117681 173113
rect 117709 173085 117744 173113
rect 117584 173051 117744 173085
rect 117584 173023 117619 173051
rect 117647 173023 117681 173051
rect 117709 173023 117744 173051
rect 117584 172989 117744 173023
rect 117584 172961 117619 172989
rect 117647 172961 117681 172989
rect 117709 172961 117744 172989
rect 117584 172944 117744 172961
rect 132944 173175 133104 173192
rect 132944 173147 132979 173175
rect 133007 173147 133041 173175
rect 133069 173147 133104 173175
rect 132944 173113 133104 173147
rect 132944 173085 132979 173113
rect 133007 173085 133041 173113
rect 133069 173085 133104 173113
rect 132944 173051 133104 173085
rect 132944 173023 132979 173051
rect 133007 173023 133041 173051
rect 133069 173023 133104 173051
rect 132944 172989 133104 173023
rect 132944 172961 132979 172989
rect 133007 172961 133041 172989
rect 133069 172961 133104 172989
rect 132944 172944 133104 172961
rect 148304 173175 148464 173192
rect 148304 173147 148339 173175
rect 148367 173147 148401 173175
rect 148429 173147 148464 173175
rect 148304 173113 148464 173147
rect 148304 173085 148339 173113
rect 148367 173085 148401 173113
rect 148429 173085 148464 173113
rect 148304 173051 148464 173085
rect 148304 173023 148339 173051
rect 148367 173023 148401 173051
rect 148429 173023 148464 173051
rect 148304 172989 148464 173023
rect 148304 172961 148339 172989
rect 148367 172961 148401 172989
rect 148429 172961 148464 172989
rect 148304 172944 148464 172961
rect 163664 173175 163824 173192
rect 163664 173147 163699 173175
rect 163727 173147 163761 173175
rect 163789 173147 163824 173175
rect 163664 173113 163824 173147
rect 163664 173085 163699 173113
rect 163727 173085 163761 173113
rect 163789 173085 163824 173113
rect 163664 173051 163824 173085
rect 163664 173023 163699 173051
rect 163727 173023 163761 173051
rect 163789 173023 163824 173051
rect 163664 172989 163824 173023
rect 163664 172961 163699 172989
rect 163727 172961 163761 172989
rect 163789 172961 163824 172989
rect 163664 172944 163824 172961
rect 179024 173175 179184 173192
rect 179024 173147 179059 173175
rect 179087 173147 179121 173175
rect 179149 173147 179184 173175
rect 179024 173113 179184 173147
rect 179024 173085 179059 173113
rect 179087 173085 179121 173113
rect 179149 173085 179184 173113
rect 179024 173051 179184 173085
rect 179024 173023 179059 173051
rect 179087 173023 179121 173051
rect 179149 173023 179184 173051
rect 179024 172989 179184 173023
rect 179024 172961 179059 172989
rect 179087 172961 179121 172989
rect 179149 172961 179184 172989
rect 179024 172944 179184 172961
rect 194384 173175 194544 173192
rect 194384 173147 194419 173175
rect 194447 173147 194481 173175
rect 194509 173147 194544 173175
rect 194384 173113 194544 173147
rect 194384 173085 194419 173113
rect 194447 173085 194481 173113
rect 194509 173085 194544 173113
rect 194384 173051 194544 173085
rect 194384 173023 194419 173051
rect 194447 173023 194481 173051
rect 194509 173023 194544 173051
rect 194384 172989 194544 173023
rect 194384 172961 194419 172989
rect 194447 172961 194481 172989
rect 194509 172961 194544 172989
rect 194384 172944 194544 172961
rect 209744 173175 209904 173192
rect 209744 173147 209779 173175
rect 209807 173147 209841 173175
rect 209869 173147 209904 173175
rect 209744 173113 209904 173147
rect 209744 173085 209779 173113
rect 209807 173085 209841 173113
rect 209869 173085 209904 173113
rect 209744 173051 209904 173085
rect 209744 173023 209779 173051
rect 209807 173023 209841 173051
rect 209869 173023 209904 173051
rect 209744 172989 209904 173023
rect 209744 172961 209779 172989
rect 209807 172961 209841 172989
rect 209869 172961 209904 172989
rect 209744 172944 209904 172961
rect 225104 173175 225264 173192
rect 225104 173147 225139 173175
rect 225167 173147 225201 173175
rect 225229 173147 225264 173175
rect 225104 173113 225264 173147
rect 225104 173085 225139 173113
rect 225167 173085 225201 173113
rect 225229 173085 225264 173113
rect 225104 173051 225264 173085
rect 225104 173023 225139 173051
rect 225167 173023 225201 173051
rect 225229 173023 225264 173051
rect 225104 172989 225264 173023
rect 225104 172961 225139 172989
rect 225167 172961 225201 172989
rect 225229 172961 225264 172989
rect 225104 172944 225264 172961
rect 240464 173175 240624 173192
rect 240464 173147 240499 173175
rect 240527 173147 240561 173175
rect 240589 173147 240624 173175
rect 240464 173113 240624 173147
rect 240464 173085 240499 173113
rect 240527 173085 240561 173113
rect 240589 173085 240624 173113
rect 240464 173051 240624 173085
rect 240464 173023 240499 173051
rect 240527 173023 240561 173051
rect 240589 173023 240624 173051
rect 240464 172989 240624 173023
rect 240464 172961 240499 172989
rect 240527 172961 240561 172989
rect 240589 172961 240624 172989
rect 240464 172944 240624 172961
rect 255824 173175 255984 173192
rect 255824 173147 255859 173175
rect 255887 173147 255921 173175
rect 255949 173147 255984 173175
rect 255824 173113 255984 173147
rect 255824 173085 255859 173113
rect 255887 173085 255921 173113
rect 255949 173085 255984 173113
rect 255824 173051 255984 173085
rect 255824 173023 255859 173051
rect 255887 173023 255921 173051
rect 255949 173023 255984 173051
rect 255824 172989 255984 173023
rect 255824 172961 255859 172989
rect 255887 172961 255921 172989
rect 255949 172961 255984 172989
rect 255824 172944 255984 172961
rect 271184 173175 271344 173192
rect 271184 173147 271219 173175
rect 271247 173147 271281 173175
rect 271309 173147 271344 173175
rect 271184 173113 271344 173147
rect 271184 173085 271219 173113
rect 271247 173085 271281 173113
rect 271309 173085 271344 173113
rect 271184 173051 271344 173085
rect 271184 173023 271219 173051
rect 271247 173023 271281 173051
rect 271309 173023 271344 173051
rect 271184 172989 271344 173023
rect 271184 172961 271219 172989
rect 271247 172961 271281 172989
rect 271309 172961 271344 172989
rect 271184 172944 271344 172961
rect 279189 173175 279499 181961
rect 279189 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 279499 173175
rect 279189 173113 279499 173147
rect 279189 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 279499 173113
rect 279189 173051 279499 173085
rect 279189 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 279499 173051
rect 279189 172989 279499 173023
rect 279189 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 279499 172989
rect 99022 88937 99050 88942
rect 99078 171514 99106 171519
rect 99078 67802 99106 171486
rect 109904 167175 110064 167192
rect 109904 167147 109939 167175
rect 109967 167147 110001 167175
rect 110029 167147 110064 167175
rect 109904 167113 110064 167147
rect 109904 167085 109939 167113
rect 109967 167085 110001 167113
rect 110029 167085 110064 167113
rect 109904 167051 110064 167085
rect 109904 167023 109939 167051
rect 109967 167023 110001 167051
rect 110029 167023 110064 167051
rect 109904 166989 110064 167023
rect 109904 166961 109939 166989
rect 109967 166961 110001 166989
rect 110029 166961 110064 166989
rect 109904 166944 110064 166961
rect 125264 167175 125424 167192
rect 125264 167147 125299 167175
rect 125327 167147 125361 167175
rect 125389 167147 125424 167175
rect 125264 167113 125424 167147
rect 125264 167085 125299 167113
rect 125327 167085 125361 167113
rect 125389 167085 125424 167113
rect 125264 167051 125424 167085
rect 125264 167023 125299 167051
rect 125327 167023 125361 167051
rect 125389 167023 125424 167051
rect 125264 166989 125424 167023
rect 125264 166961 125299 166989
rect 125327 166961 125361 166989
rect 125389 166961 125424 166989
rect 125264 166944 125424 166961
rect 140624 167175 140784 167192
rect 140624 167147 140659 167175
rect 140687 167147 140721 167175
rect 140749 167147 140784 167175
rect 140624 167113 140784 167147
rect 140624 167085 140659 167113
rect 140687 167085 140721 167113
rect 140749 167085 140784 167113
rect 140624 167051 140784 167085
rect 140624 167023 140659 167051
rect 140687 167023 140721 167051
rect 140749 167023 140784 167051
rect 140624 166989 140784 167023
rect 140624 166961 140659 166989
rect 140687 166961 140721 166989
rect 140749 166961 140784 166989
rect 140624 166944 140784 166961
rect 155984 167175 156144 167192
rect 155984 167147 156019 167175
rect 156047 167147 156081 167175
rect 156109 167147 156144 167175
rect 155984 167113 156144 167147
rect 155984 167085 156019 167113
rect 156047 167085 156081 167113
rect 156109 167085 156144 167113
rect 155984 167051 156144 167085
rect 155984 167023 156019 167051
rect 156047 167023 156081 167051
rect 156109 167023 156144 167051
rect 155984 166989 156144 167023
rect 155984 166961 156019 166989
rect 156047 166961 156081 166989
rect 156109 166961 156144 166989
rect 155984 166944 156144 166961
rect 171344 167175 171504 167192
rect 171344 167147 171379 167175
rect 171407 167147 171441 167175
rect 171469 167147 171504 167175
rect 171344 167113 171504 167147
rect 171344 167085 171379 167113
rect 171407 167085 171441 167113
rect 171469 167085 171504 167113
rect 171344 167051 171504 167085
rect 171344 167023 171379 167051
rect 171407 167023 171441 167051
rect 171469 167023 171504 167051
rect 171344 166989 171504 167023
rect 171344 166961 171379 166989
rect 171407 166961 171441 166989
rect 171469 166961 171504 166989
rect 171344 166944 171504 166961
rect 186704 167175 186864 167192
rect 186704 167147 186739 167175
rect 186767 167147 186801 167175
rect 186829 167147 186864 167175
rect 186704 167113 186864 167147
rect 186704 167085 186739 167113
rect 186767 167085 186801 167113
rect 186829 167085 186864 167113
rect 186704 167051 186864 167085
rect 186704 167023 186739 167051
rect 186767 167023 186801 167051
rect 186829 167023 186864 167051
rect 186704 166989 186864 167023
rect 186704 166961 186739 166989
rect 186767 166961 186801 166989
rect 186829 166961 186864 166989
rect 186704 166944 186864 166961
rect 202064 167175 202224 167192
rect 202064 167147 202099 167175
rect 202127 167147 202161 167175
rect 202189 167147 202224 167175
rect 202064 167113 202224 167147
rect 202064 167085 202099 167113
rect 202127 167085 202161 167113
rect 202189 167085 202224 167113
rect 202064 167051 202224 167085
rect 202064 167023 202099 167051
rect 202127 167023 202161 167051
rect 202189 167023 202224 167051
rect 202064 166989 202224 167023
rect 202064 166961 202099 166989
rect 202127 166961 202161 166989
rect 202189 166961 202224 166989
rect 202064 166944 202224 166961
rect 217424 167175 217584 167192
rect 217424 167147 217459 167175
rect 217487 167147 217521 167175
rect 217549 167147 217584 167175
rect 217424 167113 217584 167147
rect 217424 167085 217459 167113
rect 217487 167085 217521 167113
rect 217549 167085 217584 167113
rect 217424 167051 217584 167085
rect 217424 167023 217459 167051
rect 217487 167023 217521 167051
rect 217549 167023 217584 167051
rect 217424 166989 217584 167023
rect 217424 166961 217459 166989
rect 217487 166961 217521 166989
rect 217549 166961 217584 166989
rect 217424 166944 217584 166961
rect 232784 167175 232944 167192
rect 232784 167147 232819 167175
rect 232847 167147 232881 167175
rect 232909 167147 232944 167175
rect 232784 167113 232944 167147
rect 232784 167085 232819 167113
rect 232847 167085 232881 167113
rect 232909 167085 232944 167113
rect 232784 167051 232944 167085
rect 232784 167023 232819 167051
rect 232847 167023 232881 167051
rect 232909 167023 232944 167051
rect 232784 166989 232944 167023
rect 232784 166961 232819 166989
rect 232847 166961 232881 166989
rect 232909 166961 232944 166989
rect 232784 166944 232944 166961
rect 248144 167175 248304 167192
rect 248144 167147 248179 167175
rect 248207 167147 248241 167175
rect 248269 167147 248304 167175
rect 248144 167113 248304 167147
rect 248144 167085 248179 167113
rect 248207 167085 248241 167113
rect 248269 167085 248304 167113
rect 248144 167051 248304 167085
rect 248144 167023 248179 167051
rect 248207 167023 248241 167051
rect 248269 167023 248304 167051
rect 248144 166989 248304 167023
rect 248144 166961 248179 166989
rect 248207 166961 248241 166989
rect 248269 166961 248304 166989
rect 248144 166944 248304 166961
rect 263504 167175 263664 167192
rect 263504 167147 263539 167175
rect 263567 167147 263601 167175
rect 263629 167147 263664 167175
rect 263504 167113 263664 167147
rect 263504 167085 263539 167113
rect 263567 167085 263601 167113
rect 263629 167085 263664 167113
rect 263504 167051 263664 167085
rect 263504 167023 263539 167051
rect 263567 167023 263601 167051
rect 263629 167023 263664 167051
rect 263504 166989 263664 167023
rect 263504 166961 263539 166989
rect 263567 166961 263601 166989
rect 263629 166961 263664 166989
rect 263504 166944 263664 166961
rect 278864 167175 279024 167192
rect 278864 167147 278899 167175
rect 278927 167147 278961 167175
rect 278989 167147 279024 167175
rect 278864 167113 279024 167147
rect 278864 167085 278899 167113
rect 278927 167085 278961 167113
rect 278989 167085 279024 167113
rect 278864 167051 279024 167085
rect 278864 167023 278899 167051
rect 278927 167023 278961 167051
rect 278989 167023 279024 167051
rect 278864 166989 279024 167023
rect 278864 166961 278899 166989
rect 278927 166961 278961 166989
rect 278989 166961 279024 166989
rect 278864 166944 279024 166961
rect 102224 164175 102384 164192
rect 102224 164147 102259 164175
rect 102287 164147 102321 164175
rect 102349 164147 102384 164175
rect 102224 164113 102384 164147
rect 102224 164085 102259 164113
rect 102287 164085 102321 164113
rect 102349 164085 102384 164113
rect 102224 164051 102384 164085
rect 102224 164023 102259 164051
rect 102287 164023 102321 164051
rect 102349 164023 102384 164051
rect 102224 163989 102384 164023
rect 102224 163961 102259 163989
rect 102287 163961 102321 163989
rect 102349 163961 102384 163989
rect 102224 163944 102384 163961
rect 117584 164175 117744 164192
rect 117584 164147 117619 164175
rect 117647 164147 117681 164175
rect 117709 164147 117744 164175
rect 117584 164113 117744 164147
rect 117584 164085 117619 164113
rect 117647 164085 117681 164113
rect 117709 164085 117744 164113
rect 117584 164051 117744 164085
rect 117584 164023 117619 164051
rect 117647 164023 117681 164051
rect 117709 164023 117744 164051
rect 117584 163989 117744 164023
rect 117584 163961 117619 163989
rect 117647 163961 117681 163989
rect 117709 163961 117744 163989
rect 117584 163944 117744 163961
rect 132944 164175 133104 164192
rect 132944 164147 132979 164175
rect 133007 164147 133041 164175
rect 133069 164147 133104 164175
rect 132944 164113 133104 164147
rect 132944 164085 132979 164113
rect 133007 164085 133041 164113
rect 133069 164085 133104 164113
rect 132944 164051 133104 164085
rect 132944 164023 132979 164051
rect 133007 164023 133041 164051
rect 133069 164023 133104 164051
rect 132944 163989 133104 164023
rect 132944 163961 132979 163989
rect 133007 163961 133041 163989
rect 133069 163961 133104 163989
rect 132944 163944 133104 163961
rect 148304 164175 148464 164192
rect 148304 164147 148339 164175
rect 148367 164147 148401 164175
rect 148429 164147 148464 164175
rect 148304 164113 148464 164147
rect 148304 164085 148339 164113
rect 148367 164085 148401 164113
rect 148429 164085 148464 164113
rect 148304 164051 148464 164085
rect 148304 164023 148339 164051
rect 148367 164023 148401 164051
rect 148429 164023 148464 164051
rect 148304 163989 148464 164023
rect 148304 163961 148339 163989
rect 148367 163961 148401 163989
rect 148429 163961 148464 163989
rect 148304 163944 148464 163961
rect 163664 164175 163824 164192
rect 163664 164147 163699 164175
rect 163727 164147 163761 164175
rect 163789 164147 163824 164175
rect 163664 164113 163824 164147
rect 163664 164085 163699 164113
rect 163727 164085 163761 164113
rect 163789 164085 163824 164113
rect 163664 164051 163824 164085
rect 163664 164023 163699 164051
rect 163727 164023 163761 164051
rect 163789 164023 163824 164051
rect 163664 163989 163824 164023
rect 163664 163961 163699 163989
rect 163727 163961 163761 163989
rect 163789 163961 163824 163989
rect 163664 163944 163824 163961
rect 179024 164175 179184 164192
rect 179024 164147 179059 164175
rect 179087 164147 179121 164175
rect 179149 164147 179184 164175
rect 179024 164113 179184 164147
rect 179024 164085 179059 164113
rect 179087 164085 179121 164113
rect 179149 164085 179184 164113
rect 179024 164051 179184 164085
rect 179024 164023 179059 164051
rect 179087 164023 179121 164051
rect 179149 164023 179184 164051
rect 179024 163989 179184 164023
rect 179024 163961 179059 163989
rect 179087 163961 179121 163989
rect 179149 163961 179184 163989
rect 179024 163944 179184 163961
rect 194384 164175 194544 164192
rect 194384 164147 194419 164175
rect 194447 164147 194481 164175
rect 194509 164147 194544 164175
rect 194384 164113 194544 164147
rect 194384 164085 194419 164113
rect 194447 164085 194481 164113
rect 194509 164085 194544 164113
rect 194384 164051 194544 164085
rect 194384 164023 194419 164051
rect 194447 164023 194481 164051
rect 194509 164023 194544 164051
rect 194384 163989 194544 164023
rect 194384 163961 194419 163989
rect 194447 163961 194481 163989
rect 194509 163961 194544 163989
rect 194384 163944 194544 163961
rect 209744 164175 209904 164192
rect 209744 164147 209779 164175
rect 209807 164147 209841 164175
rect 209869 164147 209904 164175
rect 209744 164113 209904 164147
rect 209744 164085 209779 164113
rect 209807 164085 209841 164113
rect 209869 164085 209904 164113
rect 209744 164051 209904 164085
rect 209744 164023 209779 164051
rect 209807 164023 209841 164051
rect 209869 164023 209904 164051
rect 209744 163989 209904 164023
rect 209744 163961 209779 163989
rect 209807 163961 209841 163989
rect 209869 163961 209904 163989
rect 209744 163944 209904 163961
rect 225104 164175 225264 164192
rect 225104 164147 225139 164175
rect 225167 164147 225201 164175
rect 225229 164147 225264 164175
rect 225104 164113 225264 164147
rect 225104 164085 225139 164113
rect 225167 164085 225201 164113
rect 225229 164085 225264 164113
rect 225104 164051 225264 164085
rect 225104 164023 225139 164051
rect 225167 164023 225201 164051
rect 225229 164023 225264 164051
rect 225104 163989 225264 164023
rect 225104 163961 225139 163989
rect 225167 163961 225201 163989
rect 225229 163961 225264 163989
rect 225104 163944 225264 163961
rect 240464 164175 240624 164192
rect 240464 164147 240499 164175
rect 240527 164147 240561 164175
rect 240589 164147 240624 164175
rect 240464 164113 240624 164147
rect 240464 164085 240499 164113
rect 240527 164085 240561 164113
rect 240589 164085 240624 164113
rect 240464 164051 240624 164085
rect 240464 164023 240499 164051
rect 240527 164023 240561 164051
rect 240589 164023 240624 164051
rect 240464 163989 240624 164023
rect 240464 163961 240499 163989
rect 240527 163961 240561 163989
rect 240589 163961 240624 163989
rect 240464 163944 240624 163961
rect 255824 164175 255984 164192
rect 255824 164147 255859 164175
rect 255887 164147 255921 164175
rect 255949 164147 255984 164175
rect 255824 164113 255984 164147
rect 255824 164085 255859 164113
rect 255887 164085 255921 164113
rect 255949 164085 255984 164113
rect 255824 164051 255984 164085
rect 255824 164023 255859 164051
rect 255887 164023 255921 164051
rect 255949 164023 255984 164051
rect 255824 163989 255984 164023
rect 255824 163961 255859 163989
rect 255887 163961 255921 163989
rect 255949 163961 255984 163989
rect 255824 163944 255984 163961
rect 271184 164175 271344 164192
rect 271184 164147 271219 164175
rect 271247 164147 271281 164175
rect 271309 164147 271344 164175
rect 271184 164113 271344 164147
rect 271184 164085 271219 164113
rect 271247 164085 271281 164113
rect 271309 164085 271344 164113
rect 271184 164051 271344 164085
rect 271184 164023 271219 164051
rect 271247 164023 271281 164051
rect 271309 164023 271344 164051
rect 271184 163989 271344 164023
rect 271184 163961 271219 163989
rect 271247 163961 271281 163989
rect 271309 163961 271344 163989
rect 271184 163944 271344 163961
rect 279189 164175 279499 172961
rect 279189 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 279499 164175
rect 279189 164113 279499 164147
rect 279189 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 279499 164113
rect 279189 164051 279499 164085
rect 279189 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 279499 164051
rect 279189 163989 279499 164023
rect 279189 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 279499 163989
rect 109904 158175 110064 158192
rect 109904 158147 109939 158175
rect 109967 158147 110001 158175
rect 110029 158147 110064 158175
rect 109904 158113 110064 158147
rect 109904 158085 109939 158113
rect 109967 158085 110001 158113
rect 110029 158085 110064 158113
rect 109904 158051 110064 158085
rect 109904 158023 109939 158051
rect 109967 158023 110001 158051
rect 110029 158023 110064 158051
rect 109904 157989 110064 158023
rect 109904 157961 109939 157989
rect 109967 157961 110001 157989
rect 110029 157961 110064 157989
rect 109904 157944 110064 157961
rect 125264 158175 125424 158192
rect 125264 158147 125299 158175
rect 125327 158147 125361 158175
rect 125389 158147 125424 158175
rect 125264 158113 125424 158147
rect 125264 158085 125299 158113
rect 125327 158085 125361 158113
rect 125389 158085 125424 158113
rect 125264 158051 125424 158085
rect 125264 158023 125299 158051
rect 125327 158023 125361 158051
rect 125389 158023 125424 158051
rect 125264 157989 125424 158023
rect 125264 157961 125299 157989
rect 125327 157961 125361 157989
rect 125389 157961 125424 157989
rect 125264 157944 125424 157961
rect 140624 158175 140784 158192
rect 140624 158147 140659 158175
rect 140687 158147 140721 158175
rect 140749 158147 140784 158175
rect 140624 158113 140784 158147
rect 140624 158085 140659 158113
rect 140687 158085 140721 158113
rect 140749 158085 140784 158113
rect 140624 158051 140784 158085
rect 140624 158023 140659 158051
rect 140687 158023 140721 158051
rect 140749 158023 140784 158051
rect 140624 157989 140784 158023
rect 140624 157961 140659 157989
rect 140687 157961 140721 157989
rect 140749 157961 140784 157989
rect 140624 157944 140784 157961
rect 155984 158175 156144 158192
rect 155984 158147 156019 158175
rect 156047 158147 156081 158175
rect 156109 158147 156144 158175
rect 155984 158113 156144 158147
rect 155984 158085 156019 158113
rect 156047 158085 156081 158113
rect 156109 158085 156144 158113
rect 155984 158051 156144 158085
rect 155984 158023 156019 158051
rect 156047 158023 156081 158051
rect 156109 158023 156144 158051
rect 155984 157989 156144 158023
rect 155984 157961 156019 157989
rect 156047 157961 156081 157989
rect 156109 157961 156144 157989
rect 155984 157944 156144 157961
rect 171344 158175 171504 158192
rect 171344 158147 171379 158175
rect 171407 158147 171441 158175
rect 171469 158147 171504 158175
rect 171344 158113 171504 158147
rect 171344 158085 171379 158113
rect 171407 158085 171441 158113
rect 171469 158085 171504 158113
rect 171344 158051 171504 158085
rect 171344 158023 171379 158051
rect 171407 158023 171441 158051
rect 171469 158023 171504 158051
rect 171344 157989 171504 158023
rect 171344 157961 171379 157989
rect 171407 157961 171441 157989
rect 171469 157961 171504 157989
rect 171344 157944 171504 157961
rect 186704 158175 186864 158192
rect 186704 158147 186739 158175
rect 186767 158147 186801 158175
rect 186829 158147 186864 158175
rect 186704 158113 186864 158147
rect 186704 158085 186739 158113
rect 186767 158085 186801 158113
rect 186829 158085 186864 158113
rect 186704 158051 186864 158085
rect 186704 158023 186739 158051
rect 186767 158023 186801 158051
rect 186829 158023 186864 158051
rect 186704 157989 186864 158023
rect 186704 157961 186739 157989
rect 186767 157961 186801 157989
rect 186829 157961 186864 157989
rect 186704 157944 186864 157961
rect 202064 158175 202224 158192
rect 202064 158147 202099 158175
rect 202127 158147 202161 158175
rect 202189 158147 202224 158175
rect 202064 158113 202224 158147
rect 202064 158085 202099 158113
rect 202127 158085 202161 158113
rect 202189 158085 202224 158113
rect 202064 158051 202224 158085
rect 202064 158023 202099 158051
rect 202127 158023 202161 158051
rect 202189 158023 202224 158051
rect 202064 157989 202224 158023
rect 202064 157961 202099 157989
rect 202127 157961 202161 157989
rect 202189 157961 202224 157989
rect 202064 157944 202224 157961
rect 217424 158175 217584 158192
rect 217424 158147 217459 158175
rect 217487 158147 217521 158175
rect 217549 158147 217584 158175
rect 217424 158113 217584 158147
rect 217424 158085 217459 158113
rect 217487 158085 217521 158113
rect 217549 158085 217584 158113
rect 217424 158051 217584 158085
rect 217424 158023 217459 158051
rect 217487 158023 217521 158051
rect 217549 158023 217584 158051
rect 217424 157989 217584 158023
rect 217424 157961 217459 157989
rect 217487 157961 217521 157989
rect 217549 157961 217584 157989
rect 217424 157944 217584 157961
rect 232784 158175 232944 158192
rect 232784 158147 232819 158175
rect 232847 158147 232881 158175
rect 232909 158147 232944 158175
rect 232784 158113 232944 158147
rect 232784 158085 232819 158113
rect 232847 158085 232881 158113
rect 232909 158085 232944 158113
rect 232784 158051 232944 158085
rect 232784 158023 232819 158051
rect 232847 158023 232881 158051
rect 232909 158023 232944 158051
rect 232784 157989 232944 158023
rect 232784 157961 232819 157989
rect 232847 157961 232881 157989
rect 232909 157961 232944 157989
rect 232784 157944 232944 157961
rect 248144 158175 248304 158192
rect 248144 158147 248179 158175
rect 248207 158147 248241 158175
rect 248269 158147 248304 158175
rect 248144 158113 248304 158147
rect 248144 158085 248179 158113
rect 248207 158085 248241 158113
rect 248269 158085 248304 158113
rect 248144 158051 248304 158085
rect 248144 158023 248179 158051
rect 248207 158023 248241 158051
rect 248269 158023 248304 158051
rect 248144 157989 248304 158023
rect 248144 157961 248179 157989
rect 248207 157961 248241 157989
rect 248269 157961 248304 157989
rect 248144 157944 248304 157961
rect 263504 158175 263664 158192
rect 263504 158147 263539 158175
rect 263567 158147 263601 158175
rect 263629 158147 263664 158175
rect 263504 158113 263664 158147
rect 263504 158085 263539 158113
rect 263567 158085 263601 158113
rect 263629 158085 263664 158113
rect 263504 158051 263664 158085
rect 263504 158023 263539 158051
rect 263567 158023 263601 158051
rect 263629 158023 263664 158051
rect 263504 157989 263664 158023
rect 263504 157961 263539 157989
rect 263567 157961 263601 157989
rect 263629 157961 263664 157989
rect 263504 157944 263664 157961
rect 278864 158175 279024 158192
rect 278864 158147 278899 158175
rect 278927 158147 278961 158175
rect 278989 158147 279024 158175
rect 278864 158113 279024 158147
rect 278864 158085 278899 158113
rect 278927 158085 278961 158113
rect 278989 158085 279024 158113
rect 278864 158051 279024 158085
rect 278864 158023 278899 158051
rect 278927 158023 278961 158051
rect 278989 158023 279024 158051
rect 278864 157989 279024 158023
rect 278864 157961 278899 157989
rect 278927 157961 278961 157989
rect 278989 157961 279024 157989
rect 278864 157944 279024 157961
rect 102224 155175 102384 155192
rect 102224 155147 102259 155175
rect 102287 155147 102321 155175
rect 102349 155147 102384 155175
rect 102224 155113 102384 155147
rect 102224 155085 102259 155113
rect 102287 155085 102321 155113
rect 102349 155085 102384 155113
rect 102224 155051 102384 155085
rect 102224 155023 102259 155051
rect 102287 155023 102321 155051
rect 102349 155023 102384 155051
rect 102224 154989 102384 155023
rect 102224 154961 102259 154989
rect 102287 154961 102321 154989
rect 102349 154961 102384 154989
rect 102224 154944 102384 154961
rect 117584 155175 117744 155192
rect 117584 155147 117619 155175
rect 117647 155147 117681 155175
rect 117709 155147 117744 155175
rect 117584 155113 117744 155147
rect 117584 155085 117619 155113
rect 117647 155085 117681 155113
rect 117709 155085 117744 155113
rect 117584 155051 117744 155085
rect 117584 155023 117619 155051
rect 117647 155023 117681 155051
rect 117709 155023 117744 155051
rect 117584 154989 117744 155023
rect 117584 154961 117619 154989
rect 117647 154961 117681 154989
rect 117709 154961 117744 154989
rect 117584 154944 117744 154961
rect 132944 155175 133104 155192
rect 132944 155147 132979 155175
rect 133007 155147 133041 155175
rect 133069 155147 133104 155175
rect 132944 155113 133104 155147
rect 132944 155085 132979 155113
rect 133007 155085 133041 155113
rect 133069 155085 133104 155113
rect 132944 155051 133104 155085
rect 132944 155023 132979 155051
rect 133007 155023 133041 155051
rect 133069 155023 133104 155051
rect 132944 154989 133104 155023
rect 132944 154961 132979 154989
rect 133007 154961 133041 154989
rect 133069 154961 133104 154989
rect 132944 154944 133104 154961
rect 148304 155175 148464 155192
rect 148304 155147 148339 155175
rect 148367 155147 148401 155175
rect 148429 155147 148464 155175
rect 148304 155113 148464 155147
rect 148304 155085 148339 155113
rect 148367 155085 148401 155113
rect 148429 155085 148464 155113
rect 148304 155051 148464 155085
rect 148304 155023 148339 155051
rect 148367 155023 148401 155051
rect 148429 155023 148464 155051
rect 148304 154989 148464 155023
rect 148304 154961 148339 154989
rect 148367 154961 148401 154989
rect 148429 154961 148464 154989
rect 148304 154944 148464 154961
rect 163664 155175 163824 155192
rect 163664 155147 163699 155175
rect 163727 155147 163761 155175
rect 163789 155147 163824 155175
rect 163664 155113 163824 155147
rect 163664 155085 163699 155113
rect 163727 155085 163761 155113
rect 163789 155085 163824 155113
rect 163664 155051 163824 155085
rect 163664 155023 163699 155051
rect 163727 155023 163761 155051
rect 163789 155023 163824 155051
rect 163664 154989 163824 155023
rect 163664 154961 163699 154989
rect 163727 154961 163761 154989
rect 163789 154961 163824 154989
rect 163664 154944 163824 154961
rect 179024 155175 179184 155192
rect 179024 155147 179059 155175
rect 179087 155147 179121 155175
rect 179149 155147 179184 155175
rect 179024 155113 179184 155147
rect 179024 155085 179059 155113
rect 179087 155085 179121 155113
rect 179149 155085 179184 155113
rect 179024 155051 179184 155085
rect 179024 155023 179059 155051
rect 179087 155023 179121 155051
rect 179149 155023 179184 155051
rect 179024 154989 179184 155023
rect 179024 154961 179059 154989
rect 179087 154961 179121 154989
rect 179149 154961 179184 154989
rect 179024 154944 179184 154961
rect 194384 155175 194544 155192
rect 194384 155147 194419 155175
rect 194447 155147 194481 155175
rect 194509 155147 194544 155175
rect 194384 155113 194544 155147
rect 194384 155085 194419 155113
rect 194447 155085 194481 155113
rect 194509 155085 194544 155113
rect 194384 155051 194544 155085
rect 194384 155023 194419 155051
rect 194447 155023 194481 155051
rect 194509 155023 194544 155051
rect 194384 154989 194544 155023
rect 194384 154961 194419 154989
rect 194447 154961 194481 154989
rect 194509 154961 194544 154989
rect 194384 154944 194544 154961
rect 209744 155175 209904 155192
rect 209744 155147 209779 155175
rect 209807 155147 209841 155175
rect 209869 155147 209904 155175
rect 209744 155113 209904 155147
rect 209744 155085 209779 155113
rect 209807 155085 209841 155113
rect 209869 155085 209904 155113
rect 209744 155051 209904 155085
rect 209744 155023 209779 155051
rect 209807 155023 209841 155051
rect 209869 155023 209904 155051
rect 209744 154989 209904 155023
rect 209744 154961 209779 154989
rect 209807 154961 209841 154989
rect 209869 154961 209904 154989
rect 209744 154944 209904 154961
rect 225104 155175 225264 155192
rect 225104 155147 225139 155175
rect 225167 155147 225201 155175
rect 225229 155147 225264 155175
rect 225104 155113 225264 155147
rect 225104 155085 225139 155113
rect 225167 155085 225201 155113
rect 225229 155085 225264 155113
rect 225104 155051 225264 155085
rect 225104 155023 225139 155051
rect 225167 155023 225201 155051
rect 225229 155023 225264 155051
rect 225104 154989 225264 155023
rect 225104 154961 225139 154989
rect 225167 154961 225201 154989
rect 225229 154961 225264 154989
rect 225104 154944 225264 154961
rect 240464 155175 240624 155192
rect 240464 155147 240499 155175
rect 240527 155147 240561 155175
rect 240589 155147 240624 155175
rect 240464 155113 240624 155147
rect 240464 155085 240499 155113
rect 240527 155085 240561 155113
rect 240589 155085 240624 155113
rect 240464 155051 240624 155085
rect 240464 155023 240499 155051
rect 240527 155023 240561 155051
rect 240589 155023 240624 155051
rect 240464 154989 240624 155023
rect 240464 154961 240499 154989
rect 240527 154961 240561 154989
rect 240589 154961 240624 154989
rect 240464 154944 240624 154961
rect 255824 155175 255984 155192
rect 255824 155147 255859 155175
rect 255887 155147 255921 155175
rect 255949 155147 255984 155175
rect 255824 155113 255984 155147
rect 255824 155085 255859 155113
rect 255887 155085 255921 155113
rect 255949 155085 255984 155113
rect 255824 155051 255984 155085
rect 255824 155023 255859 155051
rect 255887 155023 255921 155051
rect 255949 155023 255984 155051
rect 255824 154989 255984 155023
rect 255824 154961 255859 154989
rect 255887 154961 255921 154989
rect 255949 154961 255984 154989
rect 255824 154944 255984 154961
rect 271184 155175 271344 155192
rect 271184 155147 271219 155175
rect 271247 155147 271281 155175
rect 271309 155147 271344 155175
rect 271184 155113 271344 155147
rect 271184 155085 271219 155113
rect 271247 155085 271281 155113
rect 271309 155085 271344 155113
rect 271184 155051 271344 155085
rect 271184 155023 271219 155051
rect 271247 155023 271281 155051
rect 271309 155023 271344 155051
rect 271184 154989 271344 155023
rect 271184 154961 271219 154989
rect 271247 154961 271281 154989
rect 271309 154961 271344 154989
rect 271184 154944 271344 154961
rect 279189 155175 279499 163961
rect 279189 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 279499 155175
rect 279189 155113 279499 155147
rect 279189 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 279499 155113
rect 279189 155051 279499 155085
rect 279189 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 279499 155051
rect 279189 154989 279499 155023
rect 279189 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 279499 154989
rect 109904 149175 110064 149192
rect 109904 149147 109939 149175
rect 109967 149147 110001 149175
rect 110029 149147 110064 149175
rect 109904 149113 110064 149147
rect 109904 149085 109939 149113
rect 109967 149085 110001 149113
rect 110029 149085 110064 149113
rect 109904 149051 110064 149085
rect 109904 149023 109939 149051
rect 109967 149023 110001 149051
rect 110029 149023 110064 149051
rect 109904 148989 110064 149023
rect 109904 148961 109939 148989
rect 109967 148961 110001 148989
rect 110029 148961 110064 148989
rect 109904 148944 110064 148961
rect 125264 149175 125424 149192
rect 125264 149147 125299 149175
rect 125327 149147 125361 149175
rect 125389 149147 125424 149175
rect 125264 149113 125424 149147
rect 125264 149085 125299 149113
rect 125327 149085 125361 149113
rect 125389 149085 125424 149113
rect 125264 149051 125424 149085
rect 125264 149023 125299 149051
rect 125327 149023 125361 149051
rect 125389 149023 125424 149051
rect 125264 148989 125424 149023
rect 125264 148961 125299 148989
rect 125327 148961 125361 148989
rect 125389 148961 125424 148989
rect 125264 148944 125424 148961
rect 140624 149175 140784 149192
rect 140624 149147 140659 149175
rect 140687 149147 140721 149175
rect 140749 149147 140784 149175
rect 140624 149113 140784 149147
rect 140624 149085 140659 149113
rect 140687 149085 140721 149113
rect 140749 149085 140784 149113
rect 140624 149051 140784 149085
rect 140624 149023 140659 149051
rect 140687 149023 140721 149051
rect 140749 149023 140784 149051
rect 140624 148989 140784 149023
rect 140624 148961 140659 148989
rect 140687 148961 140721 148989
rect 140749 148961 140784 148989
rect 140624 148944 140784 148961
rect 155984 149175 156144 149192
rect 155984 149147 156019 149175
rect 156047 149147 156081 149175
rect 156109 149147 156144 149175
rect 155984 149113 156144 149147
rect 155984 149085 156019 149113
rect 156047 149085 156081 149113
rect 156109 149085 156144 149113
rect 155984 149051 156144 149085
rect 155984 149023 156019 149051
rect 156047 149023 156081 149051
rect 156109 149023 156144 149051
rect 155984 148989 156144 149023
rect 155984 148961 156019 148989
rect 156047 148961 156081 148989
rect 156109 148961 156144 148989
rect 155984 148944 156144 148961
rect 171344 149175 171504 149192
rect 171344 149147 171379 149175
rect 171407 149147 171441 149175
rect 171469 149147 171504 149175
rect 171344 149113 171504 149147
rect 171344 149085 171379 149113
rect 171407 149085 171441 149113
rect 171469 149085 171504 149113
rect 171344 149051 171504 149085
rect 171344 149023 171379 149051
rect 171407 149023 171441 149051
rect 171469 149023 171504 149051
rect 171344 148989 171504 149023
rect 171344 148961 171379 148989
rect 171407 148961 171441 148989
rect 171469 148961 171504 148989
rect 171344 148944 171504 148961
rect 186704 149175 186864 149192
rect 186704 149147 186739 149175
rect 186767 149147 186801 149175
rect 186829 149147 186864 149175
rect 186704 149113 186864 149147
rect 186704 149085 186739 149113
rect 186767 149085 186801 149113
rect 186829 149085 186864 149113
rect 186704 149051 186864 149085
rect 186704 149023 186739 149051
rect 186767 149023 186801 149051
rect 186829 149023 186864 149051
rect 186704 148989 186864 149023
rect 186704 148961 186739 148989
rect 186767 148961 186801 148989
rect 186829 148961 186864 148989
rect 186704 148944 186864 148961
rect 202064 149175 202224 149192
rect 202064 149147 202099 149175
rect 202127 149147 202161 149175
rect 202189 149147 202224 149175
rect 202064 149113 202224 149147
rect 202064 149085 202099 149113
rect 202127 149085 202161 149113
rect 202189 149085 202224 149113
rect 202064 149051 202224 149085
rect 202064 149023 202099 149051
rect 202127 149023 202161 149051
rect 202189 149023 202224 149051
rect 202064 148989 202224 149023
rect 202064 148961 202099 148989
rect 202127 148961 202161 148989
rect 202189 148961 202224 148989
rect 202064 148944 202224 148961
rect 217424 149175 217584 149192
rect 217424 149147 217459 149175
rect 217487 149147 217521 149175
rect 217549 149147 217584 149175
rect 217424 149113 217584 149147
rect 217424 149085 217459 149113
rect 217487 149085 217521 149113
rect 217549 149085 217584 149113
rect 217424 149051 217584 149085
rect 217424 149023 217459 149051
rect 217487 149023 217521 149051
rect 217549 149023 217584 149051
rect 217424 148989 217584 149023
rect 217424 148961 217459 148989
rect 217487 148961 217521 148989
rect 217549 148961 217584 148989
rect 217424 148944 217584 148961
rect 232784 149175 232944 149192
rect 232784 149147 232819 149175
rect 232847 149147 232881 149175
rect 232909 149147 232944 149175
rect 232784 149113 232944 149147
rect 232784 149085 232819 149113
rect 232847 149085 232881 149113
rect 232909 149085 232944 149113
rect 232784 149051 232944 149085
rect 232784 149023 232819 149051
rect 232847 149023 232881 149051
rect 232909 149023 232944 149051
rect 232784 148989 232944 149023
rect 232784 148961 232819 148989
rect 232847 148961 232881 148989
rect 232909 148961 232944 148989
rect 232784 148944 232944 148961
rect 248144 149175 248304 149192
rect 248144 149147 248179 149175
rect 248207 149147 248241 149175
rect 248269 149147 248304 149175
rect 248144 149113 248304 149147
rect 248144 149085 248179 149113
rect 248207 149085 248241 149113
rect 248269 149085 248304 149113
rect 248144 149051 248304 149085
rect 248144 149023 248179 149051
rect 248207 149023 248241 149051
rect 248269 149023 248304 149051
rect 248144 148989 248304 149023
rect 248144 148961 248179 148989
rect 248207 148961 248241 148989
rect 248269 148961 248304 148989
rect 248144 148944 248304 148961
rect 263504 149175 263664 149192
rect 263504 149147 263539 149175
rect 263567 149147 263601 149175
rect 263629 149147 263664 149175
rect 263504 149113 263664 149147
rect 263504 149085 263539 149113
rect 263567 149085 263601 149113
rect 263629 149085 263664 149113
rect 263504 149051 263664 149085
rect 263504 149023 263539 149051
rect 263567 149023 263601 149051
rect 263629 149023 263664 149051
rect 263504 148989 263664 149023
rect 263504 148961 263539 148989
rect 263567 148961 263601 148989
rect 263629 148961 263664 148989
rect 263504 148944 263664 148961
rect 278864 149175 279024 149192
rect 278864 149147 278899 149175
rect 278927 149147 278961 149175
rect 278989 149147 279024 149175
rect 278864 149113 279024 149147
rect 278864 149085 278899 149113
rect 278927 149085 278961 149113
rect 278989 149085 279024 149113
rect 278864 149051 279024 149085
rect 278864 149023 278899 149051
rect 278927 149023 278961 149051
rect 278989 149023 279024 149051
rect 278864 148989 279024 149023
rect 278864 148961 278899 148989
rect 278927 148961 278961 148989
rect 278989 148961 279024 148989
rect 278864 148944 279024 148961
rect 102224 146175 102384 146192
rect 102224 146147 102259 146175
rect 102287 146147 102321 146175
rect 102349 146147 102384 146175
rect 102224 146113 102384 146147
rect 102224 146085 102259 146113
rect 102287 146085 102321 146113
rect 102349 146085 102384 146113
rect 102224 146051 102384 146085
rect 102224 146023 102259 146051
rect 102287 146023 102321 146051
rect 102349 146023 102384 146051
rect 102224 145989 102384 146023
rect 102224 145961 102259 145989
rect 102287 145961 102321 145989
rect 102349 145961 102384 145989
rect 102224 145944 102384 145961
rect 117584 146175 117744 146192
rect 117584 146147 117619 146175
rect 117647 146147 117681 146175
rect 117709 146147 117744 146175
rect 117584 146113 117744 146147
rect 117584 146085 117619 146113
rect 117647 146085 117681 146113
rect 117709 146085 117744 146113
rect 117584 146051 117744 146085
rect 117584 146023 117619 146051
rect 117647 146023 117681 146051
rect 117709 146023 117744 146051
rect 117584 145989 117744 146023
rect 117584 145961 117619 145989
rect 117647 145961 117681 145989
rect 117709 145961 117744 145989
rect 117584 145944 117744 145961
rect 132944 146175 133104 146192
rect 132944 146147 132979 146175
rect 133007 146147 133041 146175
rect 133069 146147 133104 146175
rect 132944 146113 133104 146147
rect 132944 146085 132979 146113
rect 133007 146085 133041 146113
rect 133069 146085 133104 146113
rect 132944 146051 133104 146085
rect 132944 146023 132979 146051
rect 133007 146023 133041 146051
rect 133069 146023 133104 146051
rect 132944 145989 133104 146023
rect 132944 145961 132979 145989
rect 133007 145961 133041 145989
rect 133069 145961 133104 145989
rect 132944 145944 133104 145961
rect 148304 146175 148464 146192
rect 148304 146147 148339 146175
rect 148367 146147 148401 146175
rect 148429 146147 148464 146175
rect 148304 146113 148464 146147
rect 148304 146085 148339 146113
rect 148367 146085 148401 146113
rect 148429 146085 148464 146113
rect 148304 146051 148464 146085
rect 148304 146023 148339 146051
rect 148367 146023 148401 146051
rect 148429 146023 148464 146051
rect 148304 145989 148464 146023
rect 148304 145961 148339 145989
rect 148367 145961 148401 145989
rect 148429 145961 148464 145989
rect 148304 145944 148464 145961
rect 163664 146175 163824 146192
rect 163664 146147 163699 146175
rect 163727 146147 163761 146175
rect 163789 146147 163824 146175
rect 163664 146113 163824 146147
rect 163664 146085 163699 146113
rect 163727 146085 163761 146113
rect 163789 146085 163824 146113
rect 163664 146051 163824 146085
rect 163664 146023 163699 146051
rect 163727 146023 163761 146051
rect 163789 146023 163824 146051
rect 163664 145989 163824 146023
rect 163664 145961 163699 145989
rect 163727 145961 163761 145989
rect 163789 145961 163824 145989
rect 163664 145944 163824 145961
rect 179024 146175 179184 146192
rect 179024 146147 179059 146175
rect 179087 146147 179121 146175
rect 179149 146147 179184 146175
rect 179024 146113 179184 146147
rect 179024 146085 179059 146113
rect 179087 146085 179121 146113
rect 179149 146085 179184 146113
rect 179024 146051 179184 146085
rect 179024 146023 179059 146051
rect 179087 146023 179121 146051
rect 179149 146023 179184 146051
rect 179024 145989 179184 146023
rect 179024 145961 179059 145989
rect 179087 145961 179121 145989
rect 179149 145961 179184 145989
rect 179024 145944 179184 145961
rect 194384 146175 194544 146192
rect 194384 146147 194419 146175
rect 194447 146147 194481 146175
rect 194509 146147 194544 146175
rect 194384 146113 194544 146147
rect 194384 146085 194419 146113
rect 194447 146085 194481 146113
rect 194509 146085 194544 146113
rect 194384 146051 194544 146085
rect 194384 146023 194419 146051
rect 194447 146023 194481 146051
rect 194509 146023 194544 146051
rect 194384 145989 194544 146023
rect 194384 145961 194419 145989
rect 194447 145961 194481 145989
rect 194509 145961 194544 145989
rect 194384 145944 194544 145961
rect 209744 146175 209904 146192
rect 209744 146147 209779 146175
rect 209807 146147 209841 146175
rect 209869 146147 209904 146175
rect 209744 146113 209904 146147
rect 209744 146085 209779 146113
rect 209807 146085 209841 146113
rect 209869 146085 209904 146113
rect 209744 146051 209904 146085
rect 209744 146023 209779 146051
rect 209807 146023 209841 146051
rect 209869 146023 209904 146051
rect 209744 145989 209904 146023
rect 209744 145961 209779 145989
rect 209807 145961 209841 145989
rect 209869 145961 209904 145989
rect 209744 145944 209904 145961
rect 225104 146175 225264 146192
rect 225104 146147 225139 146175
rect 225167 146147 225201 146175
rect 225229 146147 225264 146175
rect 225104 146113 225264 146147
rect 225104 146085 225139 146113
rect 225167 146085 225201 146113
rect 225229 146085 225264 146113
rect 225104 146051 225264 146085
rect 225104 146023 225139 146051
rect 225167 146023 225201 146051
rect 225229 146023 225264 146051
rect 225104 145989 225264 146023
rect 225104 145961 225139 145989
rect 225167 145961 225201 145989
rect 225229 145961 225264 145989
rect 225104 145944 225264 145961
rect 240464 146175 240624 146192
rect 240464 146147 240499 146175
rect 240527 146147 240561 146175
rect 240589 146147 240624 146175
rect 240464 146113 240624 146147
rect 240464 146085 240499 146113
rect 240527 146085 240561 146113
rect 240589 146085 240624 146113
rect 240464 146051 240624 146085
rect 240464 146023 240499 146051
rect 240527 146023 240561 146051
rect 240589 146023 240624 146051
rect 240464 145989 240624 146023
rect 240464 145961 240499 145989
rect 240527 145961 240561 145989
rect 240589 145961 240624 145989
rect 240464 145944 240624 145961
rect 255824 146175 255984 146192
rect 255824 146147 255859 146175
rect 255887 146147 255921 146175
rect 255949 146147 255984 146175
rect 255824 146113 255984 146147
rect 255824 146085 255859 146113
rect 255887 146085 255921 146113
rect 255949 146085 255984 146113
rect 255824 146051 255984 146085
rect 255824 146023 255859 146051
rect 255887 146023 255921 146051
rect 255949 146023 255984 146051
rect 255824 145989 255984 146023
rect 255824 145961 255859 145989
rect 255887 145961 255921 145989
rect 255949 145961 255984 145989
rect 255824 145944 255984 145961
rect 271184 146175 271344 146192
rect 271184 146147 271219 146175
rect 271247 146147 271281 146175
rect 271309 146147 271344 146175
rect 271184 146113 271344 146147
rect 271184 146085 271219 146113
rect 271247 146085 271281 146113
rect 271309 146085 271344 146113
rect 271184 146051 271344 146085
rect 271184 146023 271219 146051
rect 271247 146023 271281 146051
rect 271309 146023 271344 146051
rect 271184 145989 271344 146023
rect 271184 145961 271219 145989
rect 271247 145961 271281 145989
rect 271309 145961 271344 145989
rect 271184 145944 271344 145961
rect 279189 146175 279499 154961
rect 279189 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 279499 146175
rect 279189 146113 279499 146147
rect 279189 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 279499 146113
rect 279189 146051 279499 146085
rect 279189 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 279499 146051
rect 279189 145989 279499 146023
rect 279189 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 279499 145989
rect 109904 140175 110064 140192
rect 109904 140147 109939 140175
rect 109967 140147 110001 140175
rect 110029 140147 110064 140175
rect 109904 140113 110064 140147
rect 109904 140085 109939 140113
rect 109967 140085 110001 140113
rect 110029 140085 110064 140113
rect 109904 140051 110064 140085
rect 109904 140023 109939 140051
rect 109967 140023 110001 140051
rect 110029 140023 110064 140051
rect 109904 139989 110064 140023
rect 109904 139961 109939 139989
rect 109967 139961 110001 139989
rect 110029 139961 110064 139989
rect 109904 139944 110064 139961
rect 125264 140175 125424 140192
rect 125264 140147 125299 140175
rect 125327 140147 125361 140175
rect 125389 140147 125424 140175
rect 125264 140113 125424 140147
rect 125264 140085 125299 140113
rect 125327 140085 125361 140113
rect 125389 140085 125424 140113
rect 125264 140051 125424 140085
rect 125264 140023 125299 140051
rect 125327 140023 125361 140051
rect 125389 140023 125424 140051
rect 125264 139989 125424 140023
rect 125264 139961 125299 139989
rect 125327 139961 125361 139989
rect 125389 139961 125424 139989
rect 125264 139944 125424 139961
rect 140624 140175 140784 140192
rect 140624 140147 140659 140175
rect 140687 140147 140721 140175
rect 140749 140147 140784 140175
rect 140624 140113 140784 140147
rect 140624 140085 140659 140113
rect 140687 140085 140721 140113
rect 140749 140085 140784 140113
rect 140624 140051 140784 140085
rect 140624 140023 140659 140051
rect 140687 140023 140721 140051
rect 140749 140023 140784 140051
rect 140624 139989 140784 140023
rect 140624 139961 140659 139989
rect 140687 139961 140721 139989
rect 140749 139961 140784 139989
rect 140624 139944 140784 139961
rect 155984 140175 156144 140192
rect 155984 140147 156019 140175
rect 156047 140147 156081 140175
rect 156109 140147 156144 140175
rect 155984 140113 156144 140147
rect 155984 140085 156019 140113
rect 156047 140085 156081 140113
rect 156109 140085 156144 140113
rect 155984 140051 156144 140085
rect 155984 140023 156019 140051
rect 156047 140023 156081 140051
rect 156109 140023 156144 140051
rect 155984 139989 156144 140023
rect 155984 139961 156019 139989
rect 156047 139961 156081 139989
rect 156109 139961 156144 139989
rect 155984 139944 156144 139961
rect 171344 140175 171504 140192
rect 171344 140147 171379 140175
rect 171407 140147 171441 140175
rect 171469 140147 171504 140175
rect 171344 140113 171504 140147
rect 171344 140085 171379 140113
rect 171407 140085 171441 140113
rect 171469 140085 171504 140113
rect 171344 140051 171504 140085
rect 171344 140023 171379 140051
rect 171407 140023 171441 140051
rect 171469 140023 171504 140051
rect 171344 139989 171504 140023
rect 171344 139961 171379 139989
rect 171407 139961 171441 139989
rect 171469 139961 171504 139989
rect 171344 139944 171504 139961
rect 186704 140175 186864 140192
rect 186704 140147 186739 140175
rect 186767 140147 186801 140175
rect 186829 140147 186864 140175
rect 186704 140113 186864 140147
rect 186704 140085 186739 140113
rect 186767 140085 186801 140113
rect 186829 140085 186864 140113
rect 186704 140051 186864 140085
rect 186704 140023 186739 140051
rect 186767 140023 186801 140051
rect 186829 140023 186864 140051
rect 186704 139989 186864 140023
rect 186704 139961 186739 139989
rect 186767 139961 186801 139989
rect 186829 139961 186864 139989
rect 186704 139944 186864 139961
rect 202064 140175 202224 140192
rect 202064 140147 202099 140175
rect 202127 140147 202161 140175
rect 202189 140147 202224 140175
rect 202064 140113 202224 140147
rect 202064 140085 202099 140113
rect 202127 140085 202161 140113
rect 202189 140085 202224 140113
rect 202064 140051 202224 140085
rect 202064 140023 202099 140051
rect 202127 140023 202161 140051
rect 202189 140023 202224 140051
rect 202064 139989 202224 140023
rect 202064 139961 202099 139989
rect 202127 139961 202161 139989
rect 202189 139961 202224 139989
rect 202064 139944 202224 139961
rect 217424 140175 217584 140192
rect 217424 140147 217459 140175
rect 217487 140147 217521 140175
rect 217549 140147 217584 140175
rect 217424 140113 217584 140147
rect 217424 140085 217459 140113
rect 217487 140085 217521 140113
rect 217549 140085 217584 140113
rect 217424 140051 217584 140085
rect 217424 140023 217459 140051
rect 217487 140023 217521 140051
rect 217549 140023 217584 140051
rect 217424 139989 217584 140023
rect 217424 139961 217459 139989
rect 217487 139961 217521 139989
rect 217549 139961 217584 139989
rect 217424 139944 217584 139961
rect 232784 140175 232944 140192
rect 232784 140147 232819 140175
rect 232847 140147 232881 140175
rect 232909 140147 232944 140175
rect 232784 140113 232944 140147
rect 232784 140085 232819 140113
rect 232847 140085 232881 140113
rect 232909 140085 232944 140113
rect 232784 140051 232944 140085
rect 232784 140023 232819 140051
rect 232847 140023 232881 140051
rect 232909 140023 232944 140051
rect 232784 139989 232944 140023
rect 232784 139961 232819 139989
rect 232847 139961 232881 139989
rect 232909 139961 232944 139989
rect 232784 139944 232944 139961
rect 248144 140175 248304 140192
rect 248144 140147 248179 140175
rect 248207 140147 248241 140175
rect 248269 140147 248304 140175
rect 248144 140113 248304 140147
rect 248144 140085 248179 140113
rect 248207 140085 248241 140113
rect 248269 140085 248304 140113
rect 248144 140051 248304 140085
rect 248144 140023 248179 140051
rect 248207 140023 248241 140051
rect 248269 140023 248304 140051
rect 248144 139989 248304 140023
rect 248144 139961 248179 139989
rect 248207 139961 248241 139989
rect 248269 139961 248304 139989
rect 248144 139944 248304 139961
rect 263504 140175 263664 140192
rect 263504 140147 263539 140175
rect 263567 140147 263601 140175
rect 263629 140147 263664 140175
rect 263504 140113 263664 140147
rect 263504 140085 263539 140113
rect 263567 140085 263601 140113
rect 263629 140085 263664 140113
rect 263504 140051 263664 140085
rect 263504 140023 263539 140051
rect 263567 140023 263601 140051
rect 263629 140023 263664 140051
rect 263504 139989 263664 140023
rect 263504 139961 263539 139989
rect 263567 139961 263601 139989
rect 263629 139961 263664 139989
rect 263504 139944 263664 139961
rect 278864 140175 279024 140192
rect 278864 140147 278899 140175
rect 278927 140147 278961 140175
rect 278989 140147 279024 140175
rect 278864 140113 279024 140147
rect 278864 140085 278899 140113
rect 278927 140085 278961 140113
rect 278989 140085 279024 140113
rect 278864 140051 279024 140085
rect 278864 140023 278899 140051
rect 278927 140023 278961 140051
rect 278989 140023 279024 140051
rect 278864 139989 279024 140023
rect 278864 139961 278899 139989
rect 278927 139961 278961 139989
rect 278989 139961 279024 139989
rect 278864 139944 279024 139961
rect 102224 137175 102384 137192
rect 102224 137147 102259 137175
rect 102287 137147 102321 137175
rect 102349 137147 102384 137175
rect 102224 137113 102384 137147
rect 102224 137085 102259 137113
rect 102287 137085 102321 137113
rect 102349 137085 102384 137113
rect 102224 137051 102384 137085
rect 102224 137023 102259 137051
rect 102287 137023 102321 137051
rect 102349 137023 102384 137051
rect 102224 136989 102384 137023
rect 102224 136961 102259 136989
rect 102287 136961 102321 136989
rect 102349 136961 102384 136989
rect 102224 136944 102384 136961
rect 117584 137175 117744 137192
rect 117584 137147 117619 137175
rect 117647 137147 117681 137175
rect 117709 137147 117744 137175
rect 117584 137113 117744 137147
rect 117584 137085 117619 137113
rect 117647 137085 117681 137113
rect 117709 137085 117744 137113
rect 117584 137051 117744 137085
rect 117584 137023 117619 137051
rect 117647 137023 117681 137051
rect 117709 137023 117744 137051
rect 117584 136989 117744 137023
rect 117584 136961 117619 136989
rect 117647 136961 117681 136989
rect 117709 136961 117744 136989
rect 117584 136944 117744 136961
rect 132944 137175 133104 137192
rect 132944 137147 132979 137175
rect 133007 137147 133041 137175
rect 133069 137147 133104 137175
rect 132944 137113 133104 137147
rect 132944 137085 132979 137113
rect 133007 137085 133041 137113
rect 133069 137085 133104 137113
rect 132944 137051 133104 137085
rect 132944 137023 132979 137051
rect 133007 137023 133041 137051
rect 133069 137023 133104 137051
rect 132944 136989 133104 137023
rect 132944 136961 132979 136989
rect 133007 136961 133041 136989
rect 133069 136961 133104 136989
rect 132944 136944 133104 136961
rect 148304 137175 148464 137192
rect 148304 137147 148339 137175
rect 148367 137147 148401 137175
rect 148429 137147 148464 137175
rect 148304 137113 148464 137147
rect 148304 137085 148339 137113
rect 148367 137085 148401 137113
rect 148429 137085 148464 137113
rect 148304 137051 148464 137085
rect 148304 137023 148339 137051
rect 148367 137023 148401 137051
rect 148429 137023 148464 137051
rect 148304 136989 148464 137023
rect 148304 136961 148339 136989
rect 148367 136961 148401 136989
rect 148429 136961 148464 136989
rect 148304 136944 148464 136961
rect 163664 137175 163824 137192
rect 163664 137147 163699 137175
rect 163727 137147 163761 137175
rect 163789 137147 163824 137175
rect 163664 137113 163824 137147
rect 163664 137085 163699 137113
rect 163727 137085 163761 137113
rect 163789 137085 163824 137113
rect 163664 137051 163824 137085
rect 163664 137023 163699 137051
rect 163727 137023 163761 137051
rect 163789 137023 163824 137051
rect 163664 136989 163824 137023
rect 163664 136961 163699 136989
rect 163727 136961 163761 136989
rect 163789 136961 163824 136989
rect 163664 136944 163824 136961
rect 179024 137175 179184 137192
rect 179024 137147 179059 137175
rect 179087 137147 179121 137175
rect 179149 137147 179184 137175
rect 179024 137113 179184 137147
rect 179024 137085 179059 137113
rect 179087 137085 179121 137113
rect 179149 137085 179184 137113
rect 179024 137051 179184 137085
rect 179024 137023 179059 137051
rect 179087 137023 179121 137051
rect 179149 137023 179184 137051
rect 179024 136989 179184 137023
rect 179024 136961 179059 136989
rect 179087 136961 179121 136989
rect 179149 136961 179184 136989
rect 179024 136944 179184 136961
rect 194384 137175 194544 137192
rect 194384 137147 194419 137175
rect 194447 137147 194481 137175
rect 194509 137147 194544 137175
rect 194384 137113 194544 137147
rect 194384 137085 194419 137113
rect 194447 137085 194481 137113
rect 194509 137085 194544 137113
rect 194384 137051 194544 137085
rect 194384 137023 194419 137051
rect 194447 137023 194481 137051
rect 194509 137023 194544 137051
rect 194384 136989 194544 137023
rect 194384 136961 194419 136989
rect 194447 136961 194481 136989
rect 194509 136961 194544 136989
rect 194384 136944 194544 136961
rect 209744 137175 209904 137192
rect 209744 137147 209779 137175
rect 209807 137147 209841 137175
rect 209869 137147 209904 137175
rect 209744 137113 209904 137147
rect 209744 137085 209779 137113
rect 209807 137085 209841 137113
rect 209869 137085 209904 137113
rect 209744 137051 209904 137085
rect 209744 137023 209779 137051
rect 209807 137023 209841 137051
rect 209869 137023 209904 137051
rect 209744 136989 209904 137023
rect 209744 136961 209779 136989
rect 209807 136961 209841 136989
rect 209869 136961 209904 136989
rect 209744 136944 209904 136961
rect 225104 137175 225264 137192
rect 225104 137147 225139 137175
rect 225167 137147 225201 137175
rect 225229 137147 225264 137175
rect 225104 137113 225264 137147
rect 225104 137085 225139 137113
rect 225167 137085 225201 137113
rect 225229 137085 225264 137113
rect 225104 137051 225264 137085
rect 225104 137023 225139 137051
rect 225167 137023 225201 137051
rect 225229 137023 225264 137051
rect 225104 136989 225264 137023
rect 225104 136961 225139 136989
rect 225167 136961 225201 136989
rect 225229 136961 225264 136989
rect 225104 136944 225264 136961
rect 240464 137175 240624 137192
rect 240464 137147 240499 137175
rect 240527 137147 240561 137175
rect 240589 137147 240624 137175
rect 240464 137113 240624 137147
rect 240464 137085 240499 137113
rect 240527 137085 240561 137113
rect 240589 137085 240624 137113
rect 240464 137051 240624 137085
rect 240464 137023 240499 137051
rect 240527 137023 240561 137051
rect 240589 137023 240624 137051
rect 240464 136989 240624 137023
rect 240464 136961 240499 136989
rect 240527 136961 240561 136989
rect 240589 136961 240624 136989
rect 240464 136944 240624 136961
rect 255824 137175 255984 137192
rect 255824 137147 255859 137175
rect 255887 137147 255921 137175
rect 255949 137147 255984 137175
rect 255824 137113 255984 137147
rect 255824 137085 255859 137113
rect 255887 137085 255921 137113
rect 255949 137085 255984 137113
rect 255824 137051 255984 137085
rect 255824 137023 255859 137051
rect 255887 137023 255921 137051
rect 255949 137023 255984 137051
rect 255824 136989 255984 137023
rect 255824 136961 255859 136989
rect 255887 136961 255921 136989
rect 255949 136961 255984 136989
rect 255824 136944 255984 136961
rect 271184 137175 271344 137192
rect 271184 137147 271219 137175
rect 271247 137147 271281 137175
rect 271309 137147 271344 137175
rect 271184 137113 271344 137147
rect 271184 137085 271219 137113
rect 271247 137085 271281 137113
rect 271309 137085 271344 137113
rect 271184 137051 271344 137085
rect 271184 137023 271219 137051
rect 271247 137023 271281 137051
rect 271309 137023 271344 137051
rect 271184 136989 271344 137023
rect 271184 136961 271219 136989
rect 271247 136961 271281 136989
rect 271309 136961 271344 136989
rect 271184 136944 271344 136961
rect 279189 137175 279499 145961
rect 279189 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 279499 137175
rect 279189 137113 279499 137147
rect 279189 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 279499 137113
rect 279189 137051 279499 137085
rect 279189 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 279499 137051
rect 279189 136989 279499 137023
rect 279189 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 279499 136989
rect 109904 131175 110064 131192
rect 109904 131147 109939 131175
rect 109967 131147 110001 131175
rect 110029 131147 110064 131175
rect 109904 131113 110064 131147
rect 109904 131085 109939 131113
rect 109967 131085 110001 131113
rect 110029 131085 110064 131113
rect 109904 131051 110064 131085
rect 109904 131023 109939 131051
rect 109967 131023 110001 131051
rect 110029 131023 110064 131051
rect 109904 130989 110064 131023
rect 109904 130961 109939 130989
rect 109967 130961 110001 130989
rect 110029 130961 110064 130989
rect 109904 130944 110064 130961
rect 125264 131175 125424 131192
rect 125264 131147 125299 131175
rect 125327 131147 125361 131175
rect 125389 131147 125424 131175
rect 125264 131113 125424 131147
rect 125264 131085 125299 131113
rect 125327 131085 125361 131113
rect 125389 131085 125424 131113
rect 125264 131051 125424 131085
rect 125264 131023 125299 131051
rect 125327 131023 125361 131051
rect 125389 131023 125424 131051
rect 125264 130989 125424 131023
rect 125264 130961 125299 130989
rect 125327 130961 125361 130989
rect 125389 130961 125424 130989
rect 125264 130944 125424 130961
rect 140624 131175 140784 131192
rect 140624 131147 140659 131175
rect 140687 131147 140721 131175
rect 140749 131147 140784 131175
rect 140624 131113 140784 131147
rect 140624 131085 140659 131113
rect 140687 131085 140721 131113
rect 140749 131085 140784 131113
rect 140624 131051 140784 131085
rect 140624 131023 140659 131051
rect 140687 131023 140721 131051
rect 140749 131023 140784 131051
rect 140624 130989 140784 131023
rect 140624 130961 140659 130989
rect 140687 130961 140721 130989
rect 140749 130961 140784 130989
rect 140624 130944 140784 130961
rect 155984 131175 156144 131192
rect 155984 131147 156019 131175
rect 156047 131147 156081 131175
rect 156109 131147 156144 131175
rect 155984 131113 156144 131147
rect 155984 131085 156019 131113
rect 156047 131085 156081 131113
rect 156109 131085 156144 131113
rect 155984 131051 156144 131085
rect 155984 131023 156019 131051
rect 156047 131023 156081 131051
rect 156109 131023 156144 131051
rect 155984 130989 156144 131023
rect 155984 130961 156019 130989
rect 156047 130961 156081 130989
rect 156109 130961 156144 130989
rect 155984 130944 156144 130961
rect 171344 131175 171504 131192
rect 171344 131147 171379 131175
rect 171407 131147 171441 131175
rect 171469 131147 171504 131175
rect 171344 131113 171504 131147
rect 171344 131085 171379 131113
rect 171407 131085 171441 131113
rect 171469 131085 171504 131113
rect 171344 131051 171504 131085
rect 171344 131023 171379 131051
rect 171407 131023 171441 131051
rect 171469 131023 171504 131051
rect 171344 130989 171504 131023
rect 171344 130961 171379 130989
rect 171407 130961 171441 130989
rect 171469 130961 171504 130989
rect 171344 130944 171504 130961
rect 186704 131175 186864 131192
rect 186704 131147 186739 131175
rect 186767 131147 186801 131175
rect 186829 131147 186864 131175
rect 186704 131113 186864 131147
rect 186704 131085 186739 131113
rect 186767 131085 186801 131113
rect 186829 131085 186864 131113
rect 186704 131051 186864 131085
rect 186704 131023 186739 131051
rect 186767 131023 186801 131051
rect 186829 131023 186864 131051
rect 186704 130989 186864 131023
rect 186704 130961 186739 130989
rect 186767 130961 186801 130989
rect 186829 130961 186864 130989
rect 186704 130944 186864 130961
rect 202064 131175 202224 131192
rect 202064 131147 202099 131175
rect 202127 131147 202161 131175
rect 202189 131147 202224 131175
rect 202064 131113 202224 131147
rect 202064 131085 202099 131113
rect 202127 131085 202161 131113
rect 202189 131085 202224 131113
rect 202064 131051 202224 131085
rect 202064 131023 202099 131051
rect 202127 131023 202161 131051
rect 202189 131023 202224 131051
rect 202064 130989 202224 131023
rect 202064 130961 202099 130989
rect 202127 130961 202161 130989
rect 202189 130961 202224 130989
rect 202064 130944 202224 130961
rect 217424 131175 217584 131192
rect 217424 131147 217459 131175
rect 217487 131147 217521 131175
rect 217549 131147 217584 131175
rect 217424 131113 217584 131147
rect 217424 131085 217459 131113
rect 217487 131085 217521 131113
rect 217549 131085 217584 131113
rect 217424 131051 217584 131085
rect 217424 131023 217459 131051
rect 217487 131023 217521 131051
rect 217549 131023 217584 131051
rect 217424 130989 217584 131023
rect 217424 130961 217459 130989
rect 217487 130961 217521 130989
rect 217549 130961 217584 130989
rect 217424 130944 217584 130961
rect 232784 131175 232944 131192
rect 232784 131147 232819 131175
rect 232847 131147 232881 131175
rect 232909 131147 232944 131175
rect 232784 131113 232944 131147
rect 232784 131085 232819 131113
rect 232847 131085 232881 131113
rect 232909 131085 232944 131113
rect 232784 131051 232944 131085
rect 232784 131023 232819 131051
rect 232847 131023 232881 131051
rect 232909 131023 232944 131051
rect 232784 130989 232944 131023
rect 232784 130961 232819 130989
rect 232847 130961 232881 130989
rect 232909 130961 232944 130989
rect 232784 130944 232944 130961
rect 248144 131175 248304 131192
rect 248144 131147 248179 131175
rect 248207 131147 248241 131175
rect 248269 131147 248304 131175
rect 248144 131113 248304 131147
rect 248144 131085 248179 131113
rect 248207 131085 248241 131113
rect 248269 131085 248304 131113
rect 248144 131051 248304 131085
rect 248144 131023 248179 131051
rect 248207 131023 248241 131051
rect 248269 131023 248304 131051
rect 248144 130989 248304 131023
rect 248144 130961 248179 130989
rect 248207 130961 248241 130989
rect 248269 130961 248304 130989
rect 248144 130944 248304 130961
rect 263504 131175 263664 131192
rect 263504 131147 263539 131175
rect 263567 131147 263601 131175
rect 263629 131147 263664 131175
rect 263504 131113 263664 131147
rect 263504 131085 263539 131113
rect 263567 131085 263601 131113
rect 263629 131085 263664 131113
rect 263504 131051 263664 131085
rect 263504 131023 263539 131051
rect 263567 131023 263601 131051
rect 263629 131023 263664 131051
rect 263504 130989 263664 131023
rect 263504 130961 263539 130989
rect 263567 130961 263601 130989
rect 263629 130961 263664 130989
rect 263504 130944 263664 130961
rect 278864 131175 279024 131192
rect 278864 131147 278899 131175
rect 278927 131147 278961 131175
rect 278989 131147 279024 131175
rect 278864 131113 279024 131147
rect 278864 131085 278899 131113
rect 278927 131085 278961 131113
rect 278989 131085 279024 131113
rect 278864 131051 279024 131085
rect 278864 131023 278899 131051
rect 278927 131023 278961 131051
rect 278989 131023 279024 131051
rect 278864 130989 279024 131023
rect 278864 130961 278899 130989
rect 278927 130961 278961 130989
rect 278989 130961 279024 130989
rect 278864 130944 279024 130961
rect 102224 128175 102384 128192
rect 102224 128147 102259 128175
rect 102287 128147 102321 128175
rect 102349 128147 102384 128175
rect 102224 128113 102384 128147
rect 102224 128085 102259 128113
rect 102287 128085 102321 128113
rect 102349 128085 102384 128113
rect 102224 128051 102384 128085
rect 102224 128023 102259 128051
rect 102287 128023 102321 128051
rect 102349 128023 102384 128051
rect 102224 127989 102384 128023
rect 102224 127961 102259 127989
rect 102287 127961 102321 127989
rect 102349 127961 102384 127989
rect 102224 127944 102384 127961
rect 117584 128175 117744 128192
rect 117584 128147 117619 128175
rect 117647 128147 117681 128175
rect 117709 128147 117744 128175
rect 117584 128113 117744 128147
rect 117584 128085 117619 128113
rect 117647 128085 117681 128113
rect 117709 128085 117744 128113
rect 117584 128051 117744 128085
rect 117584 128023 117619 128051
rect 117647 128023 117681 128051
rect 117709 128023 117744 128051
rect 117584 127989 117744 128023
rect 117584 127961 117619 127989
rect 117647 127961 117681 127989
rect 117709 127961 117744 127989
rect 117584 127944 117744 127961
rect 132944 128175 133104 128192
rect 132944 128147 132979 128175
rect 133007 128147 133041 128175
rect 133069 128147 133104 128175
rect 132944 128113 133104 128147
rect 132944 128085 132979 128113
rect 133007 128085 133041 128113
rect 133069 128085 133104 128113
rect 132944 128051 133104 128085
rect 132944 128023 132979 128051
rect 133007 128023 133041 128051
rect 133069 128023 133104 128051
rect 132944 127989 133104 128023
rect 132944 127961 132979 127989
rect 133007 127961 133041 127989
rect 133069 127961 133104 127989
rect 132944 127944 133104 127961
rect 148304 128175 148464 128192
rect 148304 128147 148339 128175
rect 148367 128147 148401 128175
rect 148429 128147 148464 128175
rect 148304 128113 148464 128147
rect 148304 128085 148339 128113
rect 148367 128085 148401 128113
rect 148429 128085 148464 128113
rect 148304 128051 148464 128085
rect 148304 128023 148339 128051
rect 148367 128023 148401 128051
rect 148429 128023 148464 128051
rect 148304 127989 148464 128023
rect 148304 127961 148339 127989
rect 148367 127961 148401 127989
rect 148429 127961 148464 127989
rect 148304 127944 148464 127961
rect 163664 128175 163824 128192
rect 163664 128147 163699 128175
rect 163727 128147 163761 128175
rect 163789 128147 163824 128175
rect 163664 128113 163824 128147
rect 163664 128085 163699 128113
rect 163727 128085 163761 128113
rect 163789 128085 163824 128113
rect 163664 128051 163824 128085
rect 163664 128023 163699 128051
rect 163727 128023 163761 128051
rect 163789 128023 163824 128051
rect 163664 127989 163824 128023
rect 163664 127961 163699 127989
rect 163727 127961 163761 127989
rect 163789 127961 163824 127989
rect 163664 127944 163824 127961
rect 179024 128175 179184 128192
rect 179024 128147 179059 128175
rect 179087 128147 179121 128175
rect 179149 128147 179184 128175
rect 179024 128113 179184 128147
rect 179024 128085 179059 128113
rect 179087 128085 179121 128113
rect 179149 128085 179184 128113
rect 179024 128051 179184 128085
rect 179024 128023 179059 128051
rect 179087 128023 179121 128051
rect 179149 128023 179184 128051
rect 179024 127989 179184 128023
rect 179024 127961 179059 127989
rect 179087 127961 179121 127989
rect 179149 127961 179184 127989
rect 179024 127944 179184 127961
rect 194384 128175 194544 128192
rect 194384 128147 194419 128175
rect 194447 128147 194481 128175
rect 194509 128147 194544 128175
rect 194384 128113 194544 128147
rect 194384 128085 194419 128113
rect 194447 128085 194481 128113
rect 194509 128085 194544 128113
rect 194384 128051 194544 128085
rect 194384 128023 194419 128051
rect 194447 128023 194481 128051
rect 194509 128023 194544 128051
rect 194384 127989 194544 128023
rect 194384 127961 194419 127989
rect 194447 127961 194481 127989
rect 194509 127961 194544 127989
rect 194384 127944 194544 127961
rect 209744 128175 209904 128192
rect 209744 128147 209779 128175
rect 209807 128147 209841 128175
rect 209869 128147 209904 128175
rect 209744 128113 209904 128147
rect 209744 128085 209779 128113
rect 209807 128085 209841 128113
rect 209869 128085 209904 128113
rect 209744 128051 209904 128085
rect 209744 128023 209779 128051
rect 209807 128023 209841 128051
rect 209869 128023 209904 128051
rect 209744 127989 209904 128023
rect 209744 127961 209779 127989
rect 209807 127961 209841 127989
rect 209869 127961 209904 127989
rect 209744 127944 209904 127961
rect 225104 128175 225264 128192
rect 225104 128147 225139 128175
rect 225167 128147 225201 128175
rect 225229 128147 225264 128175
rect 225104 128113 225264 128147
rect 225104 128085 225139 128113
rect 225167 128085 225201 128113
rect 225229 128085 225264 128113
rect 225104 128051 225264 128085
rect 225104 128023 225139 128051
rect 225167 128023 225201 128051
rect 225229 128023 225264 128051
rect 225104 127989 225264 128023
rect 225104 127961 225139 127989
rect 225167 127961 225201 127989
rect 225229 127961 225264 127989
rect 225104 127944 225264 127961
rect 240464 128175 240624 128192
rect 240464 128147 240499 128175
rect 240527 128147 240561 128175
rect 240589 128147 240624 128175
rect 240464 128113 240624 128147
rect 240464 128085 240499 128113
rect 240527 128085 240561 128113
rect 240589 128085 240624 128113
rect 240464 128051 240624 128085
rect 240464 128023 240499 128051
rect 240527 128023 240561 128051
rect 240589 128023 240624 128051
rect 240464 127989 240624 128023
rect 240464 127961 240499 127989
rect 240527 127961 240561 127989
rect 240589 127961 240624 127989
rect 240464 127944 240624 127961
rect 255824 128175 255984 128192
rect 255824 128147 255859 128175
rect 255887 128147 255921 128175
rect 255949 128147 255984 128175
rect 255824 128113 255984 128147
rect 255824 128085 255859 128113
rect 255887 128085 255921 128113
rect 255949 128085 255984 128113
rect 255824 128051 255984 128085
rect 255824 128023 255859 128051
rect 255887 128023 255921 128051
rect 255949 128023 255984 128051
rect 255824 127989 255984 128023
rect 255824 127961 255859 127989
rect 255887 127961 255921 127989
rect 255949 127961 255984 127989
rect 255824 127944 255984 127961
rect 271184 128175 271344 128192
rect 271184 128147 271219 128175
rect 271247 128147 271281 128175
rect 271309 128147 271344 128175
rect 271184 128113 271344 128147
rect 271184 128085 271219 128113
rect 271247 128085 271281 128113
rect 271309 128085 271344 128113
rect 271184 128051 271344 128085
rect 271184 128023 271219 128051
rect 271247 128023 271281 128051
rect 271309 128023 271344 128051
rect 271184 127989 271344 128023
rect 271184 127961 271219 127989
rect 271247 127961 271281 127989
rect 271309 127961 271344 127989
rect 271184 127944 271344 127961
rect 279189 128175 279499 136961
rect 279189 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 279499 128175
rect 279189 128113 279499 128147
rect 279189 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 279499 128113
rect 279189 128051 279499 128085
rect 279189 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 279499 128051
rect 279189 127989 279499 128023
rect 279189 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 279499 127989
rect 109904 122175 110064 122192
rect 109904 122147 109939 122175
rect 109967 122147 110001 122175
rect 110029 122147 110064 122175
rect 109904 122113 110064 122147
rect 109904 122085 109939 122113
rect 109967 122085 110001 122113
rect 110029 122085 110064 122113
rect 109904 122051 110064 122085
rect 109904 122023 109939 122051
rect 109967 122023 110001 122051
rect 110029 122023 110064 122051
rect 109904 121989 110064 122023
rect 109904 121961 109939 121989
rect 109967 121961 110001 121989
rect 110029 121961 110064 121989
rect 109904 121944 110064 121961
rect 125264 122175 125424 122192
rect 125264 122147 125299 122175
rect 125327 122147 125361 122175
rect 125389 122147 125424 122175
rect 125264 122113 125424 122147
rect 125264 122085 125299 122113
rect 125327 122085 125361 122113
rect 125389 122085 125424 122113
rect 125264 122051 125424 122085
rect 125264 122023 125299 122051
rect 125327 122023 125361 122051
rect 125389 122023 125424 122051
rect 125264 121989 125424 122023
rect 125264 121961 125299 121989
rect 125327 121961 125361 121989
rect 125389 121961 125424 121989
rect 125264 121944 125424 121961
rect 140624 122175 140784 122192
rect 140624 122147 140659 122175
rect 140687 122147 140721 122175
rect 140749 122147 140784 122175
rect 140624 122113 140784 122147
rect 140624 122085 140659 122113
rect 140687 122085 140721 122113
rect 140749 122085 140784 122113
rect 140624 122051 140784 122085
rect 140624 122023 140659 122051
rect 140687 122023 140721 122051
rect 140749 122023 140784 122051
rect 140624 121989 140784 122023
rect 140624 121961 140659 121989
rect 140687 121961 140721 121989
rect 140749 121961 140784 121989
rect 140624 121944 140784 121961
rect 155984 122175 156144 122192
rect 155984 122147 156019 122175
rect 156047 122147 156081 122175
rect 156109 122147 156144 122175
rect 155984 122113 156144 122147
rect 155984 122085 156019 122113
rect 156047 122085 156081 122113
rect 156109 122085 156144 122113
rect 155984 122051 156144 122085
rect 155984 122023 156019 122051
rect 156047 122023 156081 122051
rect 156109 122023 156144 122051
rect 155984 121989 156144 122023
rect 155984 121961 156019 121989
rect 156047 121961 156081 121989
rect 156109 121961 156144 121989
rect 155984 121944 156144 121961
rect 171344 122175 171504 122192
rect 171344 122147 171379 122175
rect 171407 122147 171441 122175
rect 171469 122147 171504 122175
rect 171344 122113 171504 122147
rect 171344 122085 171379 122113
rect 171407 122085 171441 122113
rect 171469 122085 171504 122113
rect 171344 122051 171504 122085
rect 171344 122023 171379 122051
rect 171407 122023 171441 122051
rect 171469 122023 171504 122051
rect 171344 121989 171504 122023
rect 171344 121961 171379 121989
rect 171407 121961 171441 121989
rect 171469 121961 171504 121989
rect 171344 121944 171504 121961
rect 186704 122175 186864 122192
rect 186704 122147 186739 122175
rect 186767 122147 186801 122175
rect 186829 122147 186864 122175
rect 186704 122113 186864 122147
rect 186704 122085 186739 122113
rect 186767 122085 186801 122113
rect 186829 122085 186864 122113
rect 186704 122051 186864 122085
rect 186704 122023 186739 122051
rect 186767 122023 186801 122051
rect 186829 122023 186864 122051
rect 186704 121989 186864 122023
rect 186704 121961 186739 121989
rect 186767 121961 186801 121989
rect 186829 121961 186864 121989
rect 186704 121944 186864 121961
rect 202064 122175 202224 122192
rect 202064 122147 202099 122175
rect 202127 122147 202161 122175
rect 202189 122147 202224 122175
rect 202064 122113 202224 122147
rect 202064 122085 202099 122113
rect 202127 122085 202161 122113
rect 202189 122085 202224 122113
rect 202064 122051 202224 122085
rect 202064 122023 202099 122051
rect 202127 122023 202161 122051
rect 202189 122023 202224 122051
rect 202064 121989 202224 122023
rect 202064 121961 202099 121989
rect 202127 121961 202161 121989
rect 202189 121961 202224 121989
rect 202064 121944 202224 121961
rect 217424 122175 217584 122192
rect 217424 122147 217459 122175
rect 217487 122147 217521 122175
rect 217549 122147 217584 122175
rect 217424 122113 217584 122147
rect 217424 122085 217459 122113
rect 217487 122085 217521 122113
rect 217549 122085 217584 122113
rect 217424 122051 217584 122085
rect 217424 122023 217459 122051
rect 217487 122023 217521 122051
rect 217549 122023 217584 122051
rect 217424 121989 217584 122023
rect 217424 121961 217459 121989
rect 217487 121961 217521 121989
rect 217549 121961 217584 121989
rect 217424 121944 217584 121961
rect 232784 122175 232944 122192
rect 232784 122147 232819 122175
rect 232847 122147 232881 122175
rect 232909 122147 232944 122175
rect 232784 122113 232944 122147
rect 232784 122085 232819 122113
rect 232847 122085 232881 122113
rect 232909 122085 232944 122113
rect 232784 122051 232944 122085
rect 232784 122023 232819 122051
rect 232847 122023 232881 122051
rect 232909 122023 232944 122051
rect 232784 121989 232944 122023
rect 232784 121961 232819 121989
rect 232847 121961 232881 121989
rect 232909 121961 232944 121989
rect 232784 121944 232944 121961
rect 248144 122175 248304 122192
rect 248144 122147 248179 122175
rect 248207 122147 248241 122175
rect 248269 122147 248304 122175
rect 248144 122113 248304 122147
rect 248144 122085 248179 122113
rect 248207 122085 248241 122113
rect 248269 122085 248304 122113
rect 248144 122051 248304 122085
rect 248144 122023 248179 122051
rect 248207 122023 248241 122051
rect 248269 122023 248304 122051
rect 248144 121989 248304 122023
rect 248144 121961 248179 121989
rect 248207 121961 248241 121989
rect 248269 121961 248304 121989
rect 248144 121944 248304 121961
rect 263504 122175 263664 122192
rect 263504 122147 263539 122175
rect 263567 122147 263601 122175
rect 263629 122147 263664 122175
rect 263504 122113 263664 122147
rect 263504 122085 263539 122113
rect 263567 122085 263601 122113
rect 263629 122085 263664 122113
rect 263504 122051 263664 122085
rect 263504 122023 263539 122051
rect 263567 122023 263601 122051
rect 263629 122023 263664 122051
rect 263504 121989 263664 122023
rect 263504 121961 263539 121989
rect 263567 121961 263601 121989
rect 263629 121961 263664 121989
rect 263504 121944 263664 121961
rect 278864 122175 279024 122192
rect 278864 122147 278899 122175
rect 278927 122147 278961 122175
rect 278989 122147 279024 122175
rect 278864 122113 279024 122147
rect 278864 122085 278899 122113
rect 278927 122085 278961 122113
rect 278989 122085 279024 122113
rect 278864 122051 279024 122085
rect 278864 122023 278899 122051
rect 278927 122023 278961 122051
rect 278989 122023 279024 122051
rect 278864 121989 279024 122023
rect 278864 121961 278899 121989
rect 278927 121961 278961 121989
rect 278989 121961 279024 121989
rect 278864 121944 279024 121961
rect 102224 119175 102384 119192
rect 102224 119147 102259 119175
rect 102287 119147 102321 119175
rect 102349 119147 102384 119175
rect 102224 119113 102384 119147
rect 102224 119085 102259 119113
rect 102287 119085 102321 119113
rect 102349 119085 102384 119113
rect 102224 119051 102384 119085
rect 102224 119023 102259 119051
rect 102287 119023 102321 119051
rect 102349 119023 102384 119051
rect 102224 118989 102384 119023
rect 102224 118961 102259 118989
rect 102287 118961 102321 118989
rect 102349 118961 102384 118989
rect 102224 118944 102384 118961
rect 117584 119175 117744 119192
rect 117584 119147 117619 119175
rect 117647 119147 117681 119175
rect 117709 119147 117744 119175
rect 117584 119113 117744 119147
rect 117584 119085 117619 119113
rect 117647 119085 117681 119113
rect 117709 119085 117744 119113
rect 117584 119051 117744 119085
rect 117584 119023 117619 119051
rect 117647 119023 117681 119051
rect 117709 119023 117744 119051
rect 117584 118989 117744 119023
rect 117584 118961 117619 118989
rect 117647 118961 117681 118989
rect 117709 118961 117744 118989
rect 117584 118944 117744 118961
rect 132944 119175 133104 119192
rect 132944 119147 132979 119175
rect 133007 119147 133041 119175
rect 133069 119147 133104 119175
rect 132944 119113 133104 119147
rect 132944 119085 132979 119113
rect 133007 119085 133041 119113
rect 133069 119085 133104 119113
rect 132944 119051 133104 119085
rect 132944 119023 132979 119051
rect 133007 119023 133041 119051
rect 133069 119023 133104 119051
rect 132944 118989 133104 119023
rect 132944 118961 132979 118989
rect 133007 118961 133041 118989
rect 133069 118961 133104 118989
rect 132944 118944 133104 118961
rect 148304 119175 148464 119192
rect 148304 119147 148339 119175
rect 148367 119147 148401 119175
rect 148429 119147 148464 119175
rect 148304 119113 148464 119147
rect 148304 119085 148339 119113
rect 148367 119085 148401 119113
rect 148429 119085 148464 119113
rect 148304 119051 148464 119085
rect 148304 119023 148339 119051
rect 148367 119023 148401 119051
rect 148429 119023 148464 119051
rect 148304 118989 148464 119023
rect 148304 118961 148339 118989
rect 148367 118961 148401 118989
rect 148429 118961 148464 118989
rect 148304 118944 148464 118961
rect 163664 119175 163824 119192
rect 163664 119147 163699 119175
rect 163727 119147 163761 119175
rect 163789 119147 163824 119175
rect 163664 119113 163824 119147
rect 163664 119085 163699 119113
rect 163727 119085 163761 119113
rect 163789 119085 163824 119113
rect 163664 119051 163824 119085
rect 163664 119023 163699 119051
rect 163727 119023 163761 119051
rect 163789 119023 163824 119051
rect 163664 118989 163824 119023
rect 163664 118961 163699 118989
rect 163727 118961 163761 118989
rect 163789 118961 163824 118989
rect 163664 118944 163824 118961
rect 179024 119175 179184 119192
rect 179024 119147 179059 119175
rect 179087 119147 179121 119175
rect 179149 119147 179184 119175
rect 179024 119113 179184 119147
rect 179024 119085 179059 119113
rect 179087 119085 179121 119113
rect 179149 119085 179184 119113
rect 179024 119051 179184 119085
rect 179024 119023 179059 119051
rect 179087 119023 179121 119051
rect 179149 119023 179184 119051
rect 179024 118989 179184 119023
rect 179024 118961 179059 118989
rect 179087 118961 179121 118989
rect 179149 118961 179184 118989
rect 179024 118944 179184 118961
rect 194384 119175 194544 119192
rect 194384 119147 194419 119175
rect 194447 119147 194481 119175
rect 194509 119147 194544 119175
rect 194384 119113 194544 119147
rect 194384 119085 194419 119113
rect 194447 119085 194481 119113
rect 194509 119085 194544 119113
rect 194384 119051 194544 119085
rect 194384 119023 194419 119051
rect 194447 119023 194481 119051
rect 194509 119023 194544 119051
rect 194384 118989 194544 119023
rect 194384 118961 194419 118989
rect 194447 118961 194481 118989
rect 194509 118961 194544 118989
rect 194384 118944 194544 118961
rect 209744 119175 209904 119192
rect 209744 119147 209779 119175
rect 209807 119147 209841 119175
rect 209869 119147 209904 119175
rect 209744 119113 209904 119147
rect 209744 119085 209779 119113
rect 209807 119085 209841 119113
rect 209869 119085 209904 119113
rect 209744 119051 209904 119085
rect 209744 119023 209779 119051
rect 209807 119023 209841 119051
rect 209869 119023 209904 119051
rect 209744 118989 209904 119023
rect 209744 118961 209779 118989
rect 209807 118961 209841 118989
rect 209869 118961 209904 118989
rect 209744 118944 209904 118961
rect 225104 119175 225264 119192
rect 225104 119147 225139 119175
rect 225167 119147 225201 119175
rect 225229 119147 225264 119175
rect 225104 119113 225264 119147
rect 225104 119085 225139 119113
rect 225167 119085 225201 119113
rect 225229 119085 225264 119113
rect 225104 119051 225264 119085
rect 225104 119023 225139 119051
rect 225167 119023 225201 119051
rect 225229 119023 225264 119051
rect 225104 118989 225264 119023
rect 225104 118961 225139 118989
rect 225167 118961 225201 118989
rect 225229 118961 225264 118989
rect 225104 118944 225264 118961
rect 240464 119175 240624 119192
rect 240464 119147 240499 119175
rect 240527 119147 240561 119175
rect 240589 119147 240624 119175
rect 240464 119113 240624 119147
rect 240464 119085 240499 119113
rect 240527 119085 240561 119113
rect 240589 119085 240624 119113
rect 240464 119051 240624 119085
rect 240464 119023 240499 119051
rect 240527 119023 240561 119051
rect 240589 119023 240624 119051
rect 240464 118989 240624 119023
rect 240464 118961 240499 118989
rect 240527 118961 240561 118989
rect 240589 118961 240624 118989
rect 240464 118944 240624 118961
rect 255824 119175 255984 119192
rect 255824 119147 255859 119175
rect 255887 119147 255921 119175
rect 255949 119147 255984 119175
rect 255824 119113 255984 119147
rect 255824 119085 255859 119113
rect 255887 119085 255921 119113
rect 255949 119085 255984 119113
rect 255824 119051 255984 119085
rect 255824 119023 255859 119051
rect 255887 119023 255921 119051
rect 255949 119023 255984 119051
rect 255824 118989 255984 119023
rect 255824 118961 255859 118989
rect 255887 118961 255921 118989
rect 255949 118961 255984 118989
rect 255824 118944 255984 118961
rect 271184 119175 271344 119192
rect 271184 119147 271219 119175
rect 271247 119147 271281 119175
rect 271309 119147 271344 119175
rect 271184 119113 271344 119147
rect 271184 119085 271219 119113
rect 271247 119085 271281 119113
rect 271309 119085 271344 119113
rect 271184 119051 271344 119085
rect 271184 119023 271219 119051
rect 271247 119023 271281 119051
rect 271309 119023 271344 119051
rect 271184 118989 271344 119023
rect 271184 118961 271219 118989
rect 271247 118961 271281 118989
rect 271309 118961 271344 118989
rect 271184 118944 271344 118961
rect 279189 119175 279499 127961
rect 279189 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 279499 119175
rect 279189 119113 279499 119147
rect 279189 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 279499 119113
rect 279189 119051 279499 119085
rect 279189 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 279499 119051
rect 279189 118989 279499 119023
rect 279189 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 279499 118989
rect 109904 113175 110064 113192
rect 109904 113147 109939 113175
rect 109967 113147 110001 113175
rect 110029 113147 110064 113175
rect 109904 113113 110064 113147
rect 109904 113085 109939 113113
rect 109967 113085 110001 113113
rect 110029 113085 110064 113113
rect 109904 113051 110064 113085
rect 109904 113023 109939 113051
rect 109967 113023 110001 113051
rect 110029 113023 110064 113051
rect 109904 112989 110064 113023
rect 109904 112961 109939 112989
rect 109967 112961 110001 112989
rect 110029 112961 110064 112989
rect 109904 112944 110064 112961
rect 125264 113175 125424 113192
rect 125264 113147 125299 113175
rect 125327 113147 125361 113175
rect 125389 113147 125424 113175
rect 125264 113113 125424 113147
rect 125264 113085 125299 113113
rect 125327 113085 125361 113113
rect 125389 113085 125424 113113
rect 125264 113051 125424 113085
rect 125264 113023 125299 113051
rect 125327 113023 125361 113051
rect 125389 113023 125424 113051
rect 125264 112989 125424 113023
rect 125264 112961 125299 112989
rect 125327 112961 125361 112989
rect 125389 112961 125424 112989
rect 125264 112944 125424 112961
rect 140624 113175 140784 113192
rect 140624 113147 140659 113175
rect 140687 113147 140721 113175
rect 140749 113147 140784 113175
rect 140624 113113 140784 113147
rect 140624 113085 140659 113113
rect 140687 113085 140721 113113
rect 140749 113085 140784 113113
rect 140624 113051 140784 113085
rect 140624 113023 140659 113051
rect 140687 113023 140721 113051
rect 140749 113023 140784 113051
rect 140624 112989 140784 113023
rect 140624 112961 140659 112989
rect 140687 112961 140721 112989
rect 140749 112961 140784 112989
rect 140624 112944 140784 112961
rect 155984 113175 156144 113192
rect 155984 113147 156019 113175
rect 156047 113147 156081 113175
rect 156109 113147 156144 113175
rect 155984 113113 156144 113147
rect 155984 113085 156019 113113
rect 156047 113085 156081 113113
rect 156109 113085 156144 113113
rect 155984 113051 156144 113085
rect 155984 113023 156019 113051
rect 156047 113023 156081 113051
rect 156109 113023 156144 113051
rect 155984 112989 156144 113023
rect 155984 112961 156019 112989
rect 156047 112961 156081 112989
rect 156109 112961 156144 112989
rect 155984 112944 156144 112961
rect 171344 113175 171504 113192
rect 171344 113147 171379 113175
rect 171407 113147 171441 113175
rect 171469 113147 171504 113175
rect 171344 113113 171504 113147
rect 171344 113085 171379 113113
rect 171407 113085 171441 113113
rect 171469 113085 171504 113113
rect 171344 113051 171504 113085
rect 171344 113023 171379 113051
rect 171407 113023 171441 113051
rect 171469 113023 171504 113051
rect 171344 112989 171504 113023
rect 171344 112961 171379 112989
rect 171407 112961 171441 112989
rect 171469 112961 171504 112989
rect 171344 112944 171504 112961
rect 186704 113175 186864 113192
rect 186704 113147 186739 113175
rect 186767 113147 186801 113175
rect 186829 113147 186864 113175
rect 186704 113113 186864 113147
rect 186704 113085 186739 113113
rect 186767 113085 186801 113113
rect 186829 113085 186864 113113
rect 186704 113051 186864 113085
rect 186704 113023 186739 113051
rect 186767 113023 186801 113051
rect 186829 113023 186864 113051
rect 186704 112989 186864 113023
rect 186704 112961 186739 112989
rect 186767 112961 186801 112989
rect 186829 112961 186864 112989
rect 186704 112944 186864 112961
rect 202064 113175 202224 113192
rect 202064 113147 202099 113175
rect 202127 113147 202161 113175
rect 202189 113147 202224 113175
rect 202064 113113 202224 113147
rect 202064 113085 202099 113113
rect 202127 113085 202161 113113
rect 202189 113085 202224 113113
rect 202064 113051 202224 113085
rect 202064 113023 202099 113051
rect 202127 113023 202161 113051
rect 202189 113023 202224 113051
rect 202064 112989 202224 113023
rect 202064 112961 202099 112989
rect 202127 112961 202161 112989
rect 202189 112961 202224 112989
rect 202064 112944 202224 112961
rect 217424 113175 217584 113192
rect 217424 113147 217459 113175
rect 217487 113147 217521 113175
rect 217549 113147 217584 113175
rect 217424 113113 217584 113147
rect 217424 113085 217459 113113
rect 217487 113085 217521 113113
rect 217549 113085 217584 113113
rect 217424 113051 217584 113085
rect 217424 113023 217459 113051
rect 217487 113023 217521 113051
rect 217549 113023 217584 113051
rect 217424 112989 217584 113023
rect 217424 112961 217459 112989
rect 217487 112961 217521 112989
rect 217549 112961 217584 112989
rect 217424 112944 217584 112961
rect 232784 113175 232944 113192
rect 232784 113147 232819 113175
rect 232847 113147 232881 113175
rect 232909 113147 232944 113175
rect 232784 113113 232944 113147
rect 232784 113085 232819 113113
rect 232847 113085 232881 113113
rect 232909 113085 232944 113113
rect 232784 113051 232944 113085
rect 232784 113023 232819 113051
rect 232847 113023 232881 113051
rect 232909 113023 232944 113051
rect 232784 112989 232944 113023
rect 232784 112961 232819 112989
rect 232847 112961 232881 112989
rect 232909 112961 232944 112989
rect 232784 112944 232944 112961
rect 248144 113175 248304 113192
rect 248144 113147 248179 113175
rect 248207 113147 248241 113175
rect 248269 113147 248304 113175
rect 248144 113113 248304 113147
rect 248144 113085 248179 113113
rect 248207 113085 248241 113113
rect 248269 113085 248304 113113
rect 248144 113051 248304 113085
rect 248144 113023 248179 113051
rect 248207 113023 248241 113051
rect 248269 113023 248304 113051
rect 248144 112989 248304 113023
rect 248144 112961 248179 112989
rect 248207 112961 248241 112989
rect 248269 112961 248304 112989
rect 248144 112944 248304 112961
rect 263504 113175 263664 113192
rect 263504 113147 263539 113175
rect 263567 113147 263601 113175
rect 263629 113147 263664 113175
rect 263504 113113 263664 113147
rect 263504 113085 263539 113113
rect 263567 113085 263601 113113
rect 263629 113085 263664 113113
rect 263504 113051 263664 113085
rect 263504 113023 263539 113051
rect 263567 113023 263601 113051
rect 263629 113023 263664 113051
rect 263504 112989 263664 113023
rect 263504 112961 263539 112989
rect 263567 112961 263601 112989
rect 263629 112961 263664 112989
rect 263504 112944 263664 112961
rect 278864 113175 279024 113192
rect 278864 113147 278899 113175
rect 278927 113147 278961 113175
rect 278989 113147 279024 113175
rect 278864 113113 279024 113147
rect 278864 113085 278899 113113
rect 278927 113085 278961 113113
rect 278989 113085 279024 113113
rect 278864 113051 279024 113085
rect 278864 113023 278899 113051
rect 278927 113023 278961 113051
rect 278989 113023 279024 113051
rect 278864 112989 279024 113023
rect 278864 112961 278899 112989
rect 278927 112961 278961 112989
rect 278989 112961 279024 112989
rect 278864 112944 279024 112961
rect 102224 110175 102384 110192
rect 102224 110147 102259 110175
rect 102287 110147 102321 110175
rect 102349 110147 102384 110175
rect 102224 110113 102384 110147
rect 102224 110085 102259 110113
rect 102287 110085 102321 110113
rect 102349 110085 102384 110113
rect 102224 110051 102384 110085
rect 102224 110023 102259 110051
rect 102287 110023 102321 110051
rect 102349 110023 102384 110051
rect 102224 109989 102384 110023
rect 102224 109961 102259 109989
rect 102287 109961 102321 109989
rect 102349 109961 102384 109989
rect 102224 109944 102384 109961
rect 117584 110175 117744 110192
rect 117584 110147 117619 110175
rect 117647 110147 117681 110175
rect 117709 110147 117744 110175
rect 117584 110113 117744 110147
rect 117584 110085 117619 110113
rect 117647 110085 117681 110113
rect 117709 110085 117744 110113
rect 117584 110051 117744 110085
rect 117584 110023 117619 110051
rect 117647 110023 117681 110051
rect 117709 110023 117744 110051
rect 117584 109989 117744 110023
rect 117584 109961 117619 109989
rect 117647 109961 117681 109989
rect 117709 109961 117744 109989
rect 117584 109944 117744 109961
rect 132944 110175 133104 110192
rect 132944 110147 132979 110175
rect 133007 110147 133041 110175
rect 133069 110147 133104 110175
rect 132944 110113 133104 110147
rect 132944 110085 132979 110113
rect 133007 110085 133041 110113
rect 133069 110085 133104 110113
rect 132944 110051 133104 110085
rect 132944 110023 132979 110051
rect 133007 110023 133041 110051
rect 133069 110023 133104 110051
rect 132944 109989 133104 110023
rect 132944 109961 132979 109989
rect 133007 109961 133041 109989
rect 133069 109961 133104 109989
rect 132944 109944 133104 109961
rect 148304 110175 148464 110192
rect 148304 110147 148339 110175
rect 148367 110147 148401 110175
rect 148429 110147 148464 110175
rect 148304 110113 148464 110147
rect 148304 110085 148339 110113
rect 148367 110085 148401 110113
rect 148429 110085 148464 110113
rect 148304 110051 148464 110085
rect 148304 110023 148339 110051
rect 148367 110023 148401 110051
rect 148429 110023 148464 110051
rect 148304 109989 148464 110023
rect 148304 109961 148339 109989
rect 148367 109961 148401 109989
rect 148429 109961 148464 109989
rect 148304 109944 148464 109961
rect 163664 110175 163824 110192
rect 163664 110147 163699 110175
rect 163727 110147 163761 110175
rect 163789 110147 163824 110175
rect 163664 110113 163824 110147
rect 163664 110085 163699 110113
rect 163727 110085 163761 110113
rect 163789 110085 163824 110113
rect 163664 110051 163824 110085
rect 163664 110023 163699 110051
rect 163727 110023 163761 110051
rect 163789 110023 163824 110051
rect 163664 109989 163824 110023
rect 163664 109961 163699 109989
rect 163727 109961 163761 109989
rect 163789 109961 163824 109989
rect 163664 109944 163824 109961
rect 179024 110175 179184 110192
rect 179024 110147 179059 110175
rect 179087 110147 179121 110175
rect 179149 110147 179184 110175
rect 179024 110113 179184 110147
rect 179024 110085 179059 110113
rect 179087 110085 179121 110113
rect 179149 110085 179184 110113
rect 179024 110051 179184 110085
rect 179024 110023 179059 110051
rect 179087 110023 179121 110051
rect 179149 110023 179184 110051
rect 179024 109989 179184 110023
rect 179024 109961 179059 109989
rect 179087 109961 179121 109989
rect 179149 109961 179184 109989
rect 179024 109944 179184 109961
rect 194384 110175 194544 110192
rect 194384 110147 194419 110175
rect 194447 110147 194481 110175
rect 194509 110147 194544 110175
rect 194384 110113 194544 110147
rect 194384 110085 194419 110113
rect 194447 110085 194481 110113
rect 194509 110085 194544 110113
rect 194384 110051 194544 110085
rect 194384 110023 194419 110051
rect 194447 110023 194481 110051
rect 194509 110023 194544 110051
rect 194384 109989 194544 110023
rect 194384 109961 194419 109989
rect 194447 109961 194481 109989
rect 194509 109961 194544 109989
rect 194384 109944 194544 109961
rect 209744 110175 209904 110192
rect 209744 110147 209779 110175
rect 209807 110147 209841 110175
rect 209869 110147 209904 110175
rect 209744 110113 209904 110147
rect 209744 110085 209779 110113
rect 209807 110085 209841 110113
rect 209869 110085 209904 110113
rect 209744 110051 209904 110085
rect 209744 110023 209779 110051
rect 209807 110023 209841 110051
rect 209869 110023 209904 110051
rect 209744 109989 209904 110023
rect 209744 109961 209779 109989
rect 209807 109961 209841 109989
rect 209869 109961 209904 109989
rect 209744 109944 209904 109961
rect 225104 110175 225264 110192
rect 225104 110147 225139 110175
rect 225167 110147 225201 110175
rect 225229 110147 225264 110175
rect 225104 110113 225264 110147
rect 225104 110085 225139 110113
rect 225167 110085 225201 110113
rect 225229 110085 225264 110113
rect 225104 110051 225264 110085
rect 225104 110023 225139 110051
rect 225167 110023 225201 110051
rect 225229 110023 225264 110051
rect 225104 109989 225264 110023
rect 225104 109961 225139 109989
rect 225167 109961 225201 109989
rect 225229 109961 225264 109989
rect 225104 109944 225264 109961
rect 240464 110175 240624 110192
rect 240464 110147 240499 110175
rect 240527 110147 240561 110175
rect 240589 110147 240624 110175
rect 240464 110113 240624 110147
rect 240464 110085 240499 110113
rect 240527 110085 240561 110113
rect 240589 110085 240624 110113
rect 240464 110051 240624 110085
rect 240464 110023 240499 110051
rect 240527 110023 240561 110051
rect 240589 110023 240624 110051
rect 240464 109989 240624 110023
rect 240464 109961 240499 109989
rect 240527 109961 240561 109989
rect 240589 109961 240624 109989
rect 240464 109944 240624 109961
rect 255824 110175 255984 110192
rect 255824 110147 255859 110175
rect 255887 110147 255921 110175
rect 255949 110147 255984 110175
rect 255824 110113 255984 110147
rect 255824 110085 255859 110113
rect 255887 110085 255921 110113
rect 255949 110085 255984 110113
rect 255824 110051 255984 110085
rect 255824 110023 255859 110051
rect 255887 110023 255921 110051
rect 255949 110023 255984 110051
rect 255824 109989 255984 110023
rect 255824 109961 255859 109989
rect 255887 109961 255921 109989
rect 255949 109961 255984 109989
rect 255824 109944 255984 109961
rect 271184 110175 271344 110192
rect 271184 110147 271219 110175
rect 271247 110147 271281 110175
rect 271309 110147 271344 110175
rect 271184 110113 271344 110147
rect 271184 110085 271219 110113
rect 271247 110085 271281 110113
rect 271309 110085 271344 110113
rect 271184 110051 271344 110085
rect 271184 110023 271219 110051
rect 271247 110023 271281 110051
rect 271309 110023 271344 110051
rect 271184 109989 271344 110023
rect 271184 109961 271219 109989
rect 271247 109961 271281 109989
rect 271309 109961 271344 109989
rect 271184 109944 271344 109961
rect 279189 110175 279499 118961
rect 279189 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 279499 110175
rect 279189 110113 279499 110147
rect 279189 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 279499 110113
rect 279189 110051 279499 110085
rect 279189 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 279499 110051
rect 279189 109989 279499 110023
rect 279189 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 279499 109989
rect 109904 104175 110064 104192
rect 109904 104147 109939 104175
rect 109967 104147 110001 104175
rect 110029 104147 110064 104175
rect 109904 104113 110064 104147
rect 109904 104085 109939 104113
rect 109967 104085 110001 104113
rect 110029 104085 110064 104113
rect 109904 104051 110064 104085
rect 109904 104023 109939 104051
rect 109967 104023 110001 104051
rect 110029 104023 110064 104051
rect 109904 103989 110064 104023
rect 109904 103961 109939 103989
rect 109967 103961 110001 103989
rect 110029 103961 110064 103989
rect 109904 103944 110064 103961
rect 125264 104175 125424 104192
rect 125264 104147 125299 104175
rect 125327 104147 125361 104175
rect 125389 104147 125424 104175
rect 125264 104113 125424 104147
rect 125264 104085 125299 104113
rect 125327 104085 125361 104113
rect 125389 104085 125424 104113
rect 125264 104051 125424 104085
rect 125264 104023 125299 104051
rect 125327 104023 125361 104051
rect 125389 104023 125424 104051
rect 125264 103989 125424 104023
rect 125264 103961 125299 103989
rect 125327 103961 125361 103989
rect 125389 103961 125424 103989
rect 125264 103944 125424 103961
rect 140624 104175 140784 104192
rect 140624 104147 140659 104175
rect 140687 104147 140721 104175
rect 140749 104147 140784 104175
rect 140624 104113 140784 104147
rect 140624 104085 140659 104113
rect 140687 104085 140721 104113
rect 140749 104085 140784 104113
rect 140624 104051 140784 104085
rect 140624 104023 140659 104051
rect 140687 104023 140721 104051
rect 140749 104023 140784 104051
rect 140624 103989 140784 104023
rect 140624 103961 140659 103989
rect 140687 103961 140721 103989
rect 140749 103961 140784 103989
rect 140624 103944 140784 103961
rect 155984 104175 156144 104192
rect 155984 104147 156019 104175
rect 156047 104147 156081 104175
rect 156109 104147 156144 104175
rect 155984 104113 156144 104147
rect 155984 104085 156019 104113
rect 156047 104085 156081 104113
rect 156109 104085 156144 104113
rect 155984 104051 156144 104085
rect 155984 104023 156019 104051
rect 156047 104023 156081 104051
rect 156109 104023 156144 104051
rect 155984 103989 156144 104023
rect 155984 103961 156019 103989
rect 156047 103961 156081 103989
rect 156109 103961 156144 103989
rect 155984 103944 156144 103961
rect 171344 104175 171504 104192
rect 171344 104147 171379 104175
rect 171407 104147 171441 104175
rect 171469 104147 171504 104175
rect 171344 104113 171504 104147
rect 171344 104085 171379 104113
rect 171407 104085 171441 104113
rect 171469 104085 171504 104113
rect 171344 104051 171504 104085
rect 171344 104023 171379 104051
rect 171407 104023 171441 104051
rect 171469 104023 171504 104051
rect 171344 103989 171504 104023
rect 171344 103961 171379 103989
rect 171407 103961 171441 103989
rect 171469 103961 171504 103989
rect 171344 103944 171504 103961
rect 186704 104175 186864 104192
rect 186704 104147 186739 104175
rect 186767 104147 186801 104175
rect 186829 104147 186864 104175
rect 186704 104113 186864 104147
rect 186704 104085 186739 104113
rect 186767 104085 186801 104113
rect 186829 104085 186864 104113
rect 186704 104051 186864 104085
rect 186704 104023 186739 104051
rect 186767 104023 186801 104051
rect 186829 104023 186864 104051
rect 186704 103989 186864 104023
rect 186704 103961 186739 103989
rect 186767 103961 186801 103989
rect 186829 103961 186864 103989
rect 186704 103944 186864 103961
rect 202064 104175 202224 104192
rect 202064 104147 202099 104175
rect 202127 104147 202161 104175
rect 202189 104147 202224 104175
rect 202064 104113 202224 104147
rect 202064 104085 202099 104113
rect 202127 104085 202161 104113
rect 202189 104085 202224 104113
rect 202064 104051 202224 104085
rect 202064 104023 202099 104051
rect 202127 104023 202161 104051
rect 202189 104023 202224 104051
rect 202064 103989 202224 104023
rect 202064 103961 202099 103989
rect 202127 103961 202161 103989
rect 202189 103961 202224 103989
rect 202064 103944 202224 103961
rect 217424 104175 217584 104192
rect 217424 104147 217459 104175
rect 217487 104147 217521 104175
rect 217549 104147 217584 104175
rect 217424 104113 217584 104147
rect 217424 104085 217459 104113
rect 217487 104085 217521 104113
rect 217549 104085 217584 104113
rect 217424 104051 217584 104085
rect 217424 104023 217459 104051
rect 217487 104023 217521 104051
rect 217549 104023 217584 104051
rect 217424 103989 217584 104023
rect 217424 103961 217459 103989
rect 217487 103961 217521 103989
rect 217549 103961 217584 103989
rect 217424 103944 217584 103961
rect 232784 104175 232944 104192
rect 232784 104147 232819 104175
rect 232847 104147 232881 104175
rect 232909 104147 232944 104175
rect 232784 104113 232944 104147
rect 232784 104085 232819 104113
rect 232847 104085 232881 104113
rect 232909 104085 232944 104113
rect 232784 104051 232944 104085
rect 232784 104023 232819 104051
rect 232847 104023 232881 104051
rect 232909 104023 232944 104051
rect 232784 103989 232944 104023
rect 232784 103961 232819 103989
rect 232847 103961 232881 103989
rect 232909 103961 232944 103989
rect 232784 103944 232944 103961
rect 248144 104175 248304 104192
rect 248144 104147 248179 104175
rect 248207 104147 248241 104175
rect 248269 104147 248304 104175
rect 248144 104113 248304 104147
rect 248144 104085 248179 104113
rect 248207 104085 248241 104113
rect 248269 104085 248304 104113
rect 248144 104051 248304 104085
rect 248144 104023 248179 104051
rect 248207 104023 248241 104051
rect 248269 104023 248304 104051
rect 248144 103989 248304 104023
rect 248144 103961 248179 103989
rect 248207 103961 248241 103989
rect 248269 103961 248304 103989
rect 248144 103944 248304 103961
rect 263504 104175 263664 104192
rect 263504 104147 263539 104175
rect 263567 104147 263601 104175
rect 263629 104147 263664 104175
rect 263504 104113 263664 104147
rect 263504 104085 263539 104113
rect 263567 104085 263601 104113
rect 263629 104085 263664 104113
rect 263504 104051 263664 104085
rect 263504 104023 263539 104051
rect 263567 104023 263601 104051
rect 263629 104023 263664 104051
rect 263504 103989 263664 104023
rect 263504 103961 263539 103989
rect 263567 103961 263601 103989
rect 263629 103961 263664 103989
rect 263504 103944 263664 103961
rect 278864 104175 279024 104192
rect 278864 104147 278899 104175
rect 278927 104147 278961 104175
rect 278989 104147 279024 104175
rect 278864 104113 279024 104147
rect 278864 104085 278899 104113
rect 278927 104085 278961 104113
rect 278989 104085 279024 104113
rect 278864 104051 279024 104085
rect 278864 104023 278899 104051
rect 278927 104023 278961 104051
rect 278989 104023 279024 104051
rect 278864 103989 279024 104023
rect 278864 103961 278899 103989
rect 278927 103961 278961 103989
rect 278989 103961 279024 103989
rect 278864 103944 279024 103961
rect 279189 101175 279499 109961
rect 279189 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 279499 101175
rect 279189 101113 279499 101147
rect 279189 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 279499 101113
rect 279189 101051 279499 101085
rect 279189 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 279499 101051
rect 279189 100989 279499 101023
rect 279189 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 279499 100989
rect 99078 67769 99106 67774
rect 110229 92175 110539 100689
rect 110229 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 110539 92175
rect 110229 92113 110539 92147
rect 110229 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 110539 92113
rect 110229 92051 110539 92085
rect 110229 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 110539 92051
rect 110229 91989 110539 92023
rect 110229 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 110539 91989
rect 110229 83175 110539 91961
rect 110229 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 110539 83175
rect 110229 83113 110539 83147
rect 110229 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 110539 83113
rect 110229 83051 110539 83085
rect 110229 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 110539 83051
rect 110229 82989 110539 83023
rect 110229 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 110539 82989
rect 110229 74175 110539 82961
rect 110229 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 110539 74175
rect 110229 74113 110539 74147
rect 110229 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 110539 74113
rect 110229 74051 110539 74085
rect 110229 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 110539 74051
rect 110229 73989 110539 74023
rect 110229 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 110539 73989
rect 98854 39545 98882 39550
rect 110229 65175 110539 73961
rect 110229 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 110539 65175
rect 110229 65113 110539 65147
rect 110229 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 110539 65113
rect 110229 65051 110539 65085
rect 110229 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 110539 65051
rect 110229 64989 110539 65023
rect 110229 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 110539 64989
rect 110229 56175 110539 64961
rect 110229 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 110539 56175
rect 110229 56113 110539 56147
rect 110229 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 110539 56113
rect 110229 56051 110539 56085
rect 110229 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 110539 56051
rect 110229 55989 110539 56023
rect 110229 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 110539 55989
rect 110229 47175 110539 55961
rect 110229 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 110539 47175
rect 110229 47113 110539 47147
rect 110229 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 110539 47113
rect 110229 47051 110539 47085
rect 110229 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 110539 47051
rect 110229 46989 110539 47023
rect 110229 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 110539 46989
rect 98798 18377 98826 18382
rect 110229 38175 110539 46961
rect 110229 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 110539 38175
rect 110229 38113 110539 38147
rect 110229 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 110539 38113
rect 110229 38051 110539 38085
rect 110229 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 110539 38051
rect 110229 37989 110539 38023
rect 110229 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 110539 37989
rect 110229 29175 110539 37961
rect 110229 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 110539 29175
rect 110229 29113 110539 29147
rect 110229 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 110539 29113
rect 110229 29051 110539 29085
rect 110229 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 110539 29051
rect 110229 28989 110539 29023
rect 110229 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 110539 28989
rect 110229 20175 110539 28961
rect 110229 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 110539 20175
rect 110229 20113 110539 20147
rect 110229 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 110539 20113
rect 110229 20051 110539 20085
rect 110229 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 110539 20051
rect 110229 19989 110539 20023
rect 110229 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 110539 19989
rect 96729 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 97039 14175
rect 96729 14113 97039 14147
rect 96729 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 97039 14113
rect 96729 14051 97039 14085
rect 96729 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 97039 14051
rect 96729 13989 97039 14023
rect 96729 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 97039 13989
rect 96729 5175 97039 13961
rect 96729 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 97039 5175
rect 96729 5113 97039 5147
rect 96729 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 97039 5113
rect 96729 5051 97039 5085
rect 96729 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 97039 5051
rect 96729 4989 97039 5023
rect 96729 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 97039 4989
rect 96729 -560 97039 4961
rect 96729 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 97039 -560
rect 96729 -622 97039 -588
rect 96729 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 97039 -622
rect 96729 -684 97039 -650
rect 96729 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 97039 -684
rect 96729 -746 97039 -712
rect 96729 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 97039 -746
rect 96729 -822 97039 -774
rect 110229 11175 110539 19961
rect 110229 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 110539 11175
rect 110229 11113 110539 11147
rect 110229 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 110539 11113
rect 110229 11051 110539 11085
rect 110229 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 110539 11051
rect 110229 10989 110539 11023
rect 110229 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 110539 10989
rect 110229 2175 110539 10961
rect 110229 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 110539 2175
rect 110229 2113 110539 2147
rect 110229 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 110539 2113
rect 110229 2051 110539 2085
rect 110229 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 110539 2051
rect 110229 1989 110539 2023
rect 110229 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 110539 1989
rect 110229 -80 110539 1961
rect 110229 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 110539 -80
rect 110229 -142 110539 -108
rect 110229 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 110539 -142
rect 110229 -204 110539 -170
rect 110229 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 110539 -204
rect 110229 -266 110539 -232
rect 110229 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 110539 -266
rect 110229 -822 110539 -294
rect 112089 95175 112399 100689
rect 112089 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 112399 95175
rect 112089 95113 112399 95147
rect 112089 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 112399 95113
rect 112089 95051 112399 95085
rect 112089 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 112399 95051
rect 112089 94989 112399 95023
rect 112089 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 112399 94989
rect 112089 86175 112399 94961
rect 112089 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 112399 86175
rect 112089 86113 112399 86147
rect 112089 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 112399 86113
rect 112089 86051 112399 86085
rect 112089 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 112399 86051
rect 112089 85989 112399 86023
rect 112089 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 112399 85989
rect 112089 77175 112399 85961
rect 112089 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 112399 77175
rect 112089 77113 112399 77147
rect 112089 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 112399 77113
rect 112089 77051 112399 77085
rect 112089 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 112399 77051
rect 112089 76989 112399 77023
rect 112089 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 112399 76989
rect 112089 68175 112399 76961
rect 112089 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 112399 68175
rect 112089 68113 112399 68147
rect 112089 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 112399 68113
rect 112089 68051 112399 68085
rect 112089 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 112399 68051
rect 112089 67989 112399 68023
rect 112089 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 112399 67989
rect 112089 59175 112399 67961
rect 112089 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 112399 59175
rect 112089 59113 112399 59147
rect 112089 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 112399 59113
rect 112089 59051 112399 59085
rect 112089 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 112399 59051
rect 112089 58989 112399 59023
rect 112089 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 112399 58989
rect 112089 50175 112399 58961
rect 112089 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 112399 50175
rect 112089 50113 112399 50147
rect 112089 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 112399 50113
rect 112089 50051 112399 50085
rect 112089 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 112399 50051
rect 112089 49989 112399 50023
rect 112089 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 112399 49989
rect 112089 41175 112399 49961
rect 112089 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 112399 41175
rect 112089 41113 112399 41147
rect 112089 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 112399 41113
rect 112089 41051 112399 41085
rect 112089 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 112399 41051
rect 112089 40989 112399 41023
rect 112089 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 112399 40989
rect 112089 32175 112399 40961
rect 112089 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 112399 32175
rect 112089 32113 112399 32147
rect 112089 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 112399 32113
rect 112089 32051 112399 32085
rect 112089 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 112399 32051
rect 112089 31989 112399 32023
rect 112089 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 112399 31989
rect 112089 23175 112399 31961
rect 112089 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 112399 23175
rect 112089 23113 112399 23147
rect 112089 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 112399 23113
rect 112089 23051 112399 23085
rect 112089 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 112399 23051
rect 112089 22989 112399 23023
rect 112089 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 112399 22989
rect 112089 14175 112399 22961
rect 112089 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 112399 14175
rect 112089 14113 112399 14147
rect 112089 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 112399 14113
rect 112089 14051 112399 14085
rect 112089 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 112399 14051
rect 112089 13989 112399 14023
rect 112089 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 112399 13989
rect 112089 5175 112399 13961
rect 112089 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 112399 5175
rect 112089 5113 112399 5147
rect 112089 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 112399 5113
rect 112089 5051 112399 5085
rect 112089 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 112399 5051
rect 112089 4989 112399 5023
rect 112089 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 112399 4989
rect 112089 -560 112399 4961
rect 112089 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 112399 -560
rect 112089 -622 112399 -588
rect 112089 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 112399 -622
rect 112089 -684 112399 -650
rect 112089 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 112399 -684
rect 112089 -746 112399 -712
rect 112089 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 112399 -746
rect 112089 -822 112399 -774
rect 125589 92175 125899 100689
rect 125589 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 125899 92175
rect 125589 92113 125899 92147
rect 125589 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 125899 92113
rect 125589 92051 125899 92085
rect 125589 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 125899 92051
rect 125589 91989 125899 92023
rect 125589 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 125899 91989
rect 125589 83175 125899 91961
rect 125589 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 125899 83175
rect 125589 83113 125899 83147
rect 125589 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 125899 83113
rect 125589 83051 125899 83085
rect 125589 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 125899 83051
rect 125589 82989 125899 83023
rect 125589 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 125899 82989
rect 125589 74175 125899 82961
rect 125589 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 125899 74175
rect 125589 74113 125899 74147
rect 125589 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 125899 74113
rect 125589 74051 125899 74085
rect 125589 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 125899 74051
rect 125589 73989 125899 74023
rect 125589 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 125899 73989
rect 125589 65175 125899 73961
rect 125589 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 125899 65175
rect 125589 65113 125899 65147
rect 125589 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 125899 65113
rect 125589 65051 125899 65085
rect 125589 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 125899 65051
rect 125589 64989 125899 65023
rect 125589 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 125899 64989
rect 125589 56175 125899 64961
rect 125589 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 125899 56175
rect 125589 56113 125899 56147
rect 125589 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 125899 56113
rect 125589 56051 125899 56085
rect 125589 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 125899 56051
rect 125589 55989 125899 56023
rect 125589 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 125899 55989
rect 125589 47175 125899 55961
rect 125589 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 125899 47175
rect 125589 47113 125899 47147
rect 125589 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 125899 47113
rect 125589 47051 125899 47085
rect 125589 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 125899 47051
rect 125589 46989 125899 47023
rect 125589 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 125899 46989
rect 125589 38175 125899 46961
rect 125589 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 125899 38175
rect 125589 38113 125899 38147
rect 125589 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 125899 38113
rect 125589 38051 125899 38085
rect 125589 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 125899 38051
rect 125589 37989 125899 38023
rect 125589 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 125899 37989
rect 125589 29175 125899 37961
rect 125589 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 125899 29175
rect 125589 29113 125899 29147
rect 125589 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 125899 29113
rect 125589 29051 125899 29085
rect 125589 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 125899 29051
rect 125589 28989 125899 29023
rect 125589 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 125899 28989
rect 125589 20175 125899 28961
rect 125589 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 125899 20175
rect 125589 20113 125899 20147
rect 125589 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 125899 20113
rect 125589 20051 125899 20085
rect 125589 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 125899 20051
rect 125589 19989 125899 20023
rect 125589 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 125899 19989
rect 125589 11175 125899 19961
rect 125589 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 125899 11175
rect 125589 11113 125899 11147
rect 125589 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 125899 11113
rect 125589 11051 125899 11085
rect 125589 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 125899 11051
rect 125589 10989 125899 11023
rect 125589 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 125899 10989
rect 125589 2175 125899 10961
rect 125589 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 125899 2175
rect 125589 2113 125899 2147
rect 125589 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 125899 2113
rect 125589 2051 125899 2085
rect 125589 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 125899 2051
rect 125589 1989 125899 2023
rect 125589 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 125899 1989
rect 125589 -80 125899 1961
rect 125589 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 125899 -80
rect 125589 -142 125899 -108
rect 125589 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 125899 -142
rect 125589 -204 125899 -170
rect 125589 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 125899 -204
rect 125589 -266 125899 -232
rect 125589 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 125899 -266
rect 125589 -822 125899 -294
rect 127449 95175 127759 100689
rect 127449 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 127759 95175
rect 127449 95113 127759 95147
rect 127449 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 127759 95113
rect 127449 95051 127759 95085
rect 127449 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 127759 95051
rect 127449 94989 127759 95023
rect 127449 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 127759 94989
rect 127449 86175 127759 94961
rect 127449 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 127759 86175
rect 127449 86113 127759 86147
rect 127449 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 127759 86113
rect 127449 86051 127759 86085
rect 127449 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 127759 86051
rect 127449 85989 127759 86023
rect 127449 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 127759 85989
rect 127449 77175 127759 85961
rect 127449 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 127759 77175
rect 127449 77113 127759 77147
rect 127449 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 127759 77113
rect 127449 77051 127759 77085
rect 127449 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 127759 77051
rect 127449 76989 127759 77023
rect 127449 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 127759 76989
rect 127449 68175 127759 76961
rect 127449 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 127759 68175
rect 127449 68113 127759 68147
rect 127449 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 127759 68113
rect 127449 68051 127759 68085
rect 127449 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 127759 68051
rect 127449 67989 127759 68023
rect 127449 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 127759 67989
rect 127449 59175 127759 67961
rect 127449 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 127759 59175
rect 127449 59113 127759 59147
rect 127449 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 127759 59113
rect 127449 59051 127759 59085
rect 127449 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 127759 59051
rect 127449 58989 127759 59023
rect 127449 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 127759 58989
rect 127449 50175 127759 58961
rect 127449 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 127759 50175
rect 127449 50113 127759 50147
rect 127449 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 127759 50113
rect 127449 50051 127759 50085
rect 127449 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 127759 50051
rect 127449 49989 127759 50023
rect 127449 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 127759 49989
rect 127449 41175 127759 49961
rect 127449 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 127759 41175
rect 127449 41113 127759 41147
rect 127449 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 127759 41113
rect 127449 41051 127759 41085
rect 127449 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 127759 41051
rect 127449 40989 127759 41023
rect 127449 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 127759 40989
rect 127449 32175 127759 40961
rect 127449 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 127759 32175
rect 127449 32113 127759 32147
rect 127449 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 127759 32113
rect 127449 32051 127759 32085
rect 127449 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 127759 32051
rect 127449 31989 127759 32023
rect 127449 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 127759 31989
rect 127449 23175 127759 31961
rect 127449 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 127759 23175
rect 127449 23113 127759 23147
rect 127449 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 127759 23113
rect 127449 23051 127759 23085
rect 127449 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 127759 23051
rect 127449 22989 127759 23023
rect 127449 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 127759 22989
rect 127449 14175 127759 22961
rect 127449 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 127759 14175
rect 127449 14113 127759 14147
rect 127449 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 127759 14113
rect 127449 14051 127759 14085
rect 127449 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 127759 14051
rect 127449 13989 127759 14023
rect 127449 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 127759 13989
rect 127449 5175 127759 13961
rect 127449 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 127759 5175
rect 127449 5113 127759 5147
rect 127449 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 127759 5113
rect 127449 5051 127759 5085
rect 127449 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 127759 5051
rect 127449 4989 127759 5023
rect 127449 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 127759 4989
rect 127449 -560 127759 4961
rect 127449 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 127759 -560
rect 127449 -622 127759 -588
rect 127449 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 127759 -622
rect 127449 -684 127759 -650
rect 127449 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 127759 -684
rect 127449 -746 127759 -712
rect 127449 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 127759 -746
rect 127449 -822 127759 -774
rect 140949 92175 141259 100689
rect 140949 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 141259 92175
rect 140949 92113 141259 92147
rect 140949 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 141259 92113
rect 140949 92051 141259 92085
rect 140949 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 141259 92051
rect 140949 91989 141259 92023
rect 140949 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 141259 91989
rect 140949 83175 141259 91961
rect 140949 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 141259 83175
rect 140949 83113 141259 83147
rect 140949 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 141259 83113
rect 140949 83051 141259 83085
rect 140949 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 141259 83051
rect 140949 82989 141259 83023
rect 140949 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 141259 82989
rect 140949 74175 141259 82961
rect 140949 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 141259 74175
rect 140949 74113 141259 74147
rect 140949 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 141259 74113
rect 140949 74051 141259 74085
rect 140949 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 141259 74051
rect 140949 73989 141259 74023
rect 140949 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 141259 73989
rect 140949 65175 141259 73961
rect 140949 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 141259 65175
rect 140949 65113 141259 65147
rect 140949 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 141259 65113
rect 140949 65051 141259 65085
rect 140949 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 141259 65051
rect 140949 64989 141259 65023
rect 140949 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 141259 64989
rect 140949 56175 141259 64961
rect 140949 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 141259 56175
rect 140949 56113 141259 56147
rect 140949 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 141259 56113
rect 140949 56051 141259 56085
rect 140949 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 141259 56051
rect 140949 55989 141259 56023
rect 140949 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 141259 55989
rect 140949 47175 141259 55961
rect 140949 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 141259 47175
rect 140949 47113 141259 47147
rect 140949 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 141259 47113
rect 140949 47051 141259 47085
rect 140949 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 141259 47051
rect 140949 46989 141259 47023
rect 140949 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 141259 46989
rect 140949 38175 141259 46961
rect 140949 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 141259 38175
rect 140949 38113 141259 38147
rect 140949 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 141259 38113
rect 140949 38051 141259 38085
rect 140949 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 141259 38051
rect 140949 37989 141259 38023
rect 140949 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 141259 37989
rect 140949 29175 141259 37961
rect 140949 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 141259 29175
rect 140949 29113 141259 29147
rect 140949 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 141259 29113
rect 140949 29051 141259 29085
rect 140949 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 141259 29051
rect 140949 28989 141259 29023
rect 140949 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 141259 28989
rect 140949 20175 141259 28961
rect 140949 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 141259 20175
rect 140949 20113 141259 20147
rect 140949 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 141259 20113
rect 140949 20051 141259 20085
rect 140949 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 141259 20051
rect 140949 19989 141259 20023
rect 140949 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 141259 19989
rect 140949 11175 141259 19961
rect 140949 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 141259 11175
rect 140949 11113 141259 11147
rect 140949 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 141259 11113
rect 140949 11051 141259 11085
rect 140949 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 141259 11051
rect 140949 10989 141259 11023
rect 140949 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 141259 10989
rect 140949 2175 141259 10961
rect 140949 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 141259 2175
rect 140949 2113 141259 2147
rect 140949 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 141259 2113
rect 140949 2051 141259 2085
rect 140949 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 141259 2051
rect 140949 1989 141259 2023
rect 140949 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 141259 1989
rect 140949 -80 141259 1961
rect 140949 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 141259 -80
rect 140949 -142 141259 -108
rect 140949 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 141259 -142
rect 140949 -204 141259 -170
rect 140949 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 141259 -204
rect 140949 -266 141259 -232
rect 140949 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 141259 -266
rect 140949 -822 141259 -294
rect 142809 95175 143119 100689
rect 142809 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 143119 95175
rect 142809 95113 143119 95147
rect 142809 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 143119 95113
rect 142809 95051 143119 95085
rect 142809 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 143119 95051
rect 142809 94989 143119 95023
rect 142809 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 143119 94989
rect 142809 86175 143119 94961
rect 142809 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 143119 86175
rect 142809 86113 143119 86147
rect 142809 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 143119 86113
rect 142809 86051 143119 86085
rect 142809 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 143119 86051
rect 142809 85989 143119 86023
rect 142809 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 143119 85989
rect 142809 77175 143119 85961
rect 142809 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 143119 77175
rect 142809 77113 143119 77147
rect 142809 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 143119 77113
rect 142809 77051 143119 77085
rect 142809 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 143119 77051
rect 142809 76989 143119 77023
rect 142809 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 143119 76989
rect 142809 68175 143119 76961
rect 142809 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 143119 68175
rect 142809 68113 143119 68147
rect 142809 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 143119 68113
rect 142809 68051 143119 68085
rect 142809 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 143119 68051
rect 142809 67989 143119 68023
rect 142809 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 143119 67989
rect 142809 59175 143119 67961
rect 142809 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 143119 59175
rect 142809 59113 143119 59147
rect 142809 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 143119 59113
rect 142809 59051 143119 59085
rect 142809 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 143119 59051
rect 142809 58989 143119 59023
rect 142809 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 143119 58989
rect 142809 50175 143119 58961
rect 142809 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 143119 50175
rect 142809 50113 143119 50147
rect 142809 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 143119 50113
rect 142809 50051 143119 50085
rect 142809 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 143119 50051
rect 142809 49989 143119 50023
rect 142809 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 143119 49989
rect 142809 41175 143119 49961
rect 142809 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 143119 41175
rect 142809 41113 143119 41147
rect 142809 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 143119 41113
rect 142809 41051 143119 41085
rect 142809 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 143119 41051
rect 142809 40989 143119 41023
rect 142809 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 143119 40989
rect 142809 32175 143119 40961
rect 142809 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 143119 32175
rect 142809 32113 143119 32147
rect 142809 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 143119 32113
rect 142809 32051 143119 32085
rect 142809 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 143119 32051
rect 142809 31989 143119 32023
rect 142809 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 143119 31989
rect 142809 23175 143119 31961
rect 142809 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 143119 23175
rect 142809 23113 143119 23147
rect 142809 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 143119 23113
rect 142809 23051 143119 23085
rect 142809 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 143119 23051
rect 142809 22989 143119 23023
rect 142809 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 143119 22989
rect 142809 14175 143119 22961
rect 142809 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 143119 14175
rect 142809 14113 143119 14147
rect 142809 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 143119 14113
rect 142809 14051 143119 14085
rect 142809 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 143119 14051
rect 142809 13989 143119 14023
rect 142809 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 143119 13989
rect 142809 5175 143119 13961
rect 142809 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 143119 5175
rect 142809 5113 143119 5147
rect 142809 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 143119 5113
rect 142809 5051 143119 5085
rect 142809 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 143119 5051
rect 142809 4989 143119 5023
rect 142809 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 143119 4989
rect 142809 -560 143119 4961
rect 142809 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 143119 -560
rect 142809 -622 143119 -588
rect 142809 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 143119 -622
rect 142809 -684 143119 -650
rect 142809 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 143119 -684
rect 142809 -746 143119 -712
rect 142809 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 143119 -746
rect 142809 -822 143119 -774
rect 156309 92175 156619 100689
rect 156309 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 156619 92175
rect 156309 92113 156619 92147
rect 156309 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 156619 92113
rect 156309 92051 156619 92085
rect 156309 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 156619 92051
rect 156309 91989 156619 92023
rect 156309 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 156619 91989
rect 156309 83175 156619 91961
rect 156309 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 156619 83175
rect 156309 83113 156619 83147
rect 156309 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 156619 83113
rect 156309 83051 156619 83085
rect 156309 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 156619 83051
rect 156309 82989 156619 83023
rect 156309 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 156619 82989
rect 156309 74175 156619 82961
rect 156309 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 156619 74175
rect 156309 74113 156619 74147
rect 156309 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 156619 74113
rect 156309 74051 156619 74085
rect 156309 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 156619 74051
rect 156309 73989 156619 74023
rect 156309 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 156619 73989
rect 156309 65175 156619 73961
rect 156309 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 156619 65175
rect 156309 65113 156619 65147
rect 156309 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 156619 65113
rect 156309 65051 156619 65085
rect 156309 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 156619 65051
rect 156309 64989 156619 65023
rect 156309 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 156619 64989
rect 156309 56175 156619 64961
rect 156309 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 156619 56175
rect 156309 56113 156619 56147
rect 156309 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 156619 56113
rect 156309 56051 156619 56085
rect 156309 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 156619 56051
rect 156309 55989 156619 56023
rect 156309 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 156619 55989
rect 156309 47175 156619 55961
rect 156309 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 156619 47175
rect 156309 47113 156619 47147
rect 156309 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 156619 47113
rect 156309 47051 156619 47085
rect 156309 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 156619 47051
rect 156309 46989 156619 47023
rect 156309 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 156619 46989
rect 156309 38175 156619 46961
rect 156309 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 156619 38175
rect 156309 38113 156619 38147
rect 156309 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 156619 38113
rect 156309 38051 156619 38085
rect 156309 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 156619 38051
rect 156309 37989 156619 38023
rect 156309 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 156619 37989
rect 156309 29175 156619 37961
rect 156309 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 156619 29175
rect 156309 29113 156619 29147
rect 156309 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 156619 29113
rect 156309 29051 156619 29085
rect 156309 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 156619 29051
rect 156309 28989 156619 29023
rect 156309 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 156619 28989
rect 156309 20175 156619 28961
rect 156309 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 156619 20175
rect 156309 20113 156619 20147
rect 156309 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 156619 20113
rect 156309 20051 156619 20085
rect 156309 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 156619 20051
rect 156309 19989 156619 20023
rect 156309 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 156619 19989
rect 156309 11175 156619 19961
rect 156309 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 156619 11175
rect 156309 11113 156619 11147
rect 156309 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 156619 11113
rect 156309 11051 156619 11085
rect 156309 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 156619 11051
rect 156309 10989 156619 11023
rect 156309 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 156619 10989
rect 156309 2175 156619 10961
rect 156309 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 156619 2175
rect 156309 2113 156619 2147
rect 156309 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 156619 2113
rect 156309 2051 156619 2085
rect 156309 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 156619 2051
rect 156309 1989 156619 2023
rect 156309 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 156619 1989
rect 156309 -80 156619 1961
rect 156309 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 156619 -80
rect 156309 -142 156619 -108
rect 156309 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 156619 -142
rect 156309 -204 156619 -170
rect 156309 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 156619 -204
rect 156309 -266 156619 -232
rect 156309 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 156619 -266
rect 156309 -822 156619 -294
rect 158169 95175 158479 100689
rect 158169 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 158479 95175
rect 158169 95113 158479 95147
rect 158169 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 158479 95113
rect 158169 95051 158479 95085
rect 158169 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 158479 95051
rect 158169 94989 158479 95023
rect 158169 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 158479 94989
rect 158169 86175 158479 94961
rect 158169 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 158479 86175
rect 158169 86113 158479 86147
rect 158169 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 158479 86113
rect 158169 86051 158479 86085
rect 158169 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 158479 86051
rect 158169 85989 158479 86023
rect 158169 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 158479 85989
rect 158169 77175 158479 85961
rect 158169 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 158479 77175
rect 158169 77113 158479 77147
rect 158169 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 158479 77113
rect 158169 77051 158479 77085
rect 158169 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 158479 77051
rect 158169 76989 158479 77023
rect 158169 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 158479 76989
rect 158169 68175 158479 76961
rect 158169 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 158479 68175
rect 158169 68113 158479 68147
rect 158169 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 158479 68113
rect 158169 68051 158479 68085
rect 158169 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 158479 68051
rect 158169 67989 158479 68023
rect 158169 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 158479 67989
rect 158169 59175 158479 67961
rect 158169 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 158479 59175
rect 158169 59113 158479 59147
rect 158169 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 158479 59113
rect 158169 59051 158479 59085
rect 158169 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 158479 59051
rect 158169 58989 158479 59023
rect 158169 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 158479 58989
rect 158169 50175 158479 58961
rect 158169 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 158479 50175
rect 158169 50113 158479 50147
rect 158169 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 158479 50113
rect 158169 50051 158479 50085
rect 158169 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 158479 50051
rect 158169 49989 158479 50023
rect 158169 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 158479 49989
rect 158169 41175 158479 49961
rect 158169 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 158479 41175
rect 158169 41113 158479 41147
rect 158169 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 158479 41113
rect 158169 41051 158479 41085
rect 158169 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 158479 41051
rect 158169 40989 158479 41023
rect 158169 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 158479 40989
rect 158169 32175 158479 40961
rect 158169 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 158479 32175
rect 158169 32113 158479 32147
rect 158169 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 158479 32113
rect 158169 32051 158479 32085
rect 158169 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 158479 32051
rect 158169 31989 158479 32023
rect 158169 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 158479 31989
rect 158169 23175 158479 31961
rect 158169 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 158479 23175
rect 158169 23113 158479 23147
rect 158169 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 158479 23113
rect 158169 23051 158479 23085
rect 158169 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 158479 23051
rect 158169 22989 158479 23023
rect 158169 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 158479 22989
rect 158169 14175 158479 22961
rect 158169 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 158479 14175
rect 158169 14113 158479 14147
rect 158169 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 158479 14113
rect 158169 14051 158479 14085
rect 158169 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 158479 14051
rect 158169 13989 158479 14023
rect 158169 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 158479 13989
rect 158169 5175 158479 13961
rect 158169 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 158479 5175
rect 158169 5113 158479 5147
rect 158169 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 158479 5113
rect 158169 5051 158479 5085
rect 158169 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 158479 5051
rect 158169 4989 158479 5023
rect 158169 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 158479 4989
rect 158169 -560 158479 4961
rect 158169 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 158479 -560
rect 158169 -622 158479 -588
rect 158169 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 158479 -622
rect 158169 -684 158479 -650
rect 158169 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 158479 -684
rect 158169 -746 158479 -712
rect 158169 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 158479 -746
rect 158169 -822 158479 -774
rect 171669 92175 171979 100689
rect 171669 92147 171717 92175
rect 171745 92147 171779 92175
rect 171807 92147 171841 92175
rect 171869 92147 171903 92175
rect 171931 92147 171979 92175
rect 171669 92113 171979 92147
rect 171669 92085 171717 92113
rect 171745 92085 171779 92113
rect 171807 92085 171841 92113
rect 171869 92085 171903 92113
rect 171931 92085 171979 92113
rect 171669 92051 171979 92085
rect 171669 92023 171717 92051
rect 171745 92023 171779 92051
rect 171807 92023 171841 92051
rect 171869 92023 171903 92051
rect 171931 92023 171979 92051
rect 171669 91989 171979 92023
rect 171669 91961 171717 91989
rect 171745 91961 171779 91989
rect 171807 91961 171841 91989
rect 171869 91961 171903 91989
rect 171931 91961 171979 91989
rect 171669 83175 171979 91961
rect 171669 83147 171717 83175
rect 171745 83147 171779 83175
rect 171807 83147 171841 83175
rect 171869 83147 171903 83175
rect 171931 83147 171979 83175
rect 171669 83113 171979 83147
rect 171669 83085 171717 83113
rect 171745 83085 171779 83113
rect 171807 83085 171841 83113
rect 171869 83085 171903 83113
rect 171931 83085 171979 83113
rect 171669 83051 171979 83085
rect 171669 83023 171717 83051
rect 171745 83023 171779 83051
rect 171807 83023 171841 83051
rect 171869 83023 171903 83051
rect 171931 83023 171979 83051
rect 171669 82989 171979 83023
rect 171669 82961 171717 82989
rect 171745 82961 171779 82989
rect 171807 82961 171841 82989
rect 171869 82961 171903 82989
rect 171931 82961 171979 82989
rect 171669 74175 171979 82961
rect 171669 74147 171717 74175
rect 171745 74147 171779 74175
rect 171807 74147 171841 74175
rect 171869 74147 171903 74175
rect 171931 74147 171979 74175
rect 171669 74113 171979 74147
rect 171669 74085 171717 74113
rect 171745 74085 171779 74113
rect 171807 74085 171841 74113
rect 171869 74085 171903 74113
rect 171931 74085 171979 74113
rect 171669 74051 171979 74085
rect 171669 74023 171717 74051
rect 171745 74023 171779 74051
rect 171807 74023 171841 74051
rect 171869 74023 171903 74051
rect 171931 74023 171979 74051
rect 171669 73989 171979 74023
rect 171669 73961 171717 73989
rect 171745 73961 171779 73989
rect 171807 73961 171841 73989
rect 171869 73961 171903 73989
rect 171931 73961 171979 73989
rect 171669 65175 171979 73961
rect 171669 65147 171717 65175
rect 171745 65147 171779 65175
rect 171807 65147 171841 65175
rect 171869 65147 171903 65175
rect 171931 65147 171979 65175
rect 171669 65113 171979 65147
rect 171669 65085 171717 65113
rect 171745 65085 171779 65113
rect 171807 65085 171841 65113
rect 171869 65085 171903 65113
rect 171931 65085 171979 65113
rect 171669 65051 171979 65085
rect 171669 65023 171717 65051
rect 171745 65023 171779 65051
rect 171807 65023 171841 65051
rect 171869 65023 171903 65051
rect 171931 65023 171979 65051
rect 171669 64989 171979 65023
rect 171669 64961 171717 64989
rect 171745 64961 171779 64989
rect 171807 64961 171841 64989
rect 171869 64961 171903 64989
rect 171931 64961 171979 64989
rect 171669 56175 171979 64961
rect 171669 56147 171717 56175
rect 171745 56147 171779 56175
rect 171807 56147 171841 56175
rect 171869 56147 171903 56175
rect 171931 56147 171979 56175
rect 171669 56113 171979 56147
rect 171669 56085 171717 56113
rect 171745 56085 171779 56113
rect 171807 56085 171841 56113
rect 171869 56085 171903 56113
rect 171931 56085 171979 56113
rect 171669 56051 171979 56085
rect 171669 56023 171717 56051
rect 171745 56023 171779 56051
rect 171807 56023 171841 56051
rect 171869 56023 171903 56051
rect 171931 56023 171979 56051
rect 171669 55989 171979 56023
rect 171669 55961 171717 55989
rect 171745 55961 171779 55989
rect 171807 55961 171841 55989
rect 171869 55961 171903 55989
rect 171931 55961 171979 55989
rect 171669 47175 171979 55961
rect 171669 47147 171717 47175
rect 171745 47147 171779 47175
rect 171807 47147 171841 47175
rect 171869 47147 171903 47175
rect 171931 47147 171979 47175
rect 171669 47113 171979 47147
rect 171669 47085 171717 47113
rect 171745 47085 171779 47113
rect 171807 47085 171841 47113
rect 171869 47085 171903 47113
rect 171931 47085 171979 47113
rect 171669 47051 171979 47085
rect 171669 47023 171717 47051
rect 171745 47023 171779 47051
rect 171807 47023 171841 47051
rect 171869 47023 171903 47051
rect 171931 47023 171979 47051
rect 171669 46989 171979 47023
rect 171669 46961 171717 46989
rect 171745 46961 171779 46989
rect 171807 46961 171841 46989
rect 171869 46961 171903 46989
rect 171931 46961 171979 46989
rect 171669 38175 171979 46961
rect 171669 38147 171717 38175
rect 171745 38147 171779 38175
rect 171807 38147 171841 38175
rect 171869 38147 171903 38175
rect 171931 38147 171979 38175
rect 171669 38113 171979 38147
rect 171669 38085 171717 38113
rect 171745 38085 171779 38113
rect 171807 38085 171841 38113
rect 171869 38085 171903 38113
rect 171931 38085 171979 38113
rect 171669 38051 171979 38085
rect 171669 38023 171717 38051
rect 171745 38023 171779 38051
rect 171807 38023 171841 38051
rect 171869 38023 171903 38051
rect 171931 38023 171979 38051
rect 171669 37989 171979 38023
rect 171669 37961 171717 37989
rect 171745 37961 171779 37989
rect 171807 37961 171841 37989
rect 171869 37961 171903 37989
rect 171931 37961 171979 37989
rect 171669 29175 171979 37961
rect 171669 29147 171717 29175
rect 171745 29147 171779 29175
rect 171807 29147 171841 29175
rect 171869 29147 171903 29175
rect 171931 29147 171979 29175
rect 171669 29113 171979 29147
rect 171669 29085 171717 29113
rect 171745 29085 171779 29113
rect 171807 29085 171841 29113
rect 171869 29085 171903 29113
rect 171931 29085 171979 29113
rect 171669 29051 171979 29085
rect 171669 29023 171717 29051
rect 171745 29023 171779 29051
rect 171807 29023 171841 29051
rect 171869 29023 171903 29051
rect 171931 29023 171979 29051
rect 171669 28989 171979 29023
rect 171669 28961 171717 28989
rect 171745 28961 171779 28989
rect 171807 28961 171841 28989
rect 171869 28961 171903 28989
rect 171931 28961 171979 28989
rect 171669 20175 171979 28961
rect 171669 20147 171717 20175
rect 171745 20147 171779 20175
rect 171807 20147 171841 20175
rect 171869 20147 171903 20175
rect 171931 20147 171979 20175
rect 171669 20113 171979 20147
rect 171669 20085 171717 20113
rect 171745 20085 171779 20113
rect 171807 20085 171841 20113
rect 171869 20085 171903 20113
rect 171931 20085 171979 20113
rect 171669 20051 171979 20085
rect 171669 20023 171717 20051
rect 171745 20023 171779 20051
rect 171807 20023 171841 20051
rect 171869 20023 171903 20051
rect 171931 20023 171979 20051
rect 171669 19989 171979 20023
rect 171669 19961 171717 19989
rect 171745 19961 171779 19989
rect 171807 19961 171841 19989
rect 171869 19961 171903 19989
rect 171931 19961 171979 19989
rect 171669 11175 171979 19961
rect 171669 11147 171717 11175
rect 171745 11147 171779 11175
rect 171807 11147 171841 11175
rect 171869 11147 171903 11175
rect 171931 11147 171979 11175
rect 171669 11113 171979 11147
rect 171669 11085 171717 11113
rect 171745 11085 171779 11113
rect 171807 11085 171841 11113
rect 171869 11085 171903 11113
rect 171931 11085 171979 11113
rect 171669 11051 171979 11085
rect 171669 11023 171717 11051
rect 171745 11023 171779 11051
rect 171807 11023 171841 11051
rect 171869 11023 171903 11051
rect 171931 11023 171979 11051
rect 171669 10989 171979 11023
rect 171669 10961 171717 10989
rect 171745 10961 171779 10989
rect 171807 10961 171841 10989
rect 171869 10961 171903 10989
rect 171931 10961 171979 10989
rect 171669 2175 171979 10961
rect 171669 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 171979 2175
rect 171669 2113 171979 2147
rect 171669 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 171979 2113
rect 171669 2051 171979 2085
rect 171669 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 171979 2051
rect 171669 1989 171979 2023
rect 171669 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 171979 1989
rect 171669 -80 171979 1961
rect 171669 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 171979 -80
rect 171669 -142 171979 -108
rect 171669 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 171979 -142
rect 171669 -204 171979 -170
rect 171669 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 171979 -204
rect 171669 -266 171979 -232
rect 171669 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 171979 -266
rect 171669 -822 171979 -294
rect 173529 95175 173839 100689
rect 173529 95147 173577 95175
rect 173605 95147 173639 95175
rect 173667 95147 173701 95175
rect 173729 95147 173763 95175
rect 173791 95147 173839 95175
rect 173529 95113 173839 95147
rect 173529 95085 173577 95113
rect 173605 95085 173639 95113
rect 173667 95085 173701 95113
rect 173729 95085 173763 95113
rect 173791 95085 173839 95113
rect 173529 95051 173839 95085
rect 173529 95023 173577 95051
rect 173605 95023 173639 95051
rect 173667 95023 173701 95051
rect 173729 95023 173763 95051
rect 173791 95023 173839 95051
rect 173529 94989 173839 95023
rect 173529 94961 173577 94989
rect 173605 94961 173639 94989
rect 173667 94961 173701 94989
rect 173729 94961 173763 94989
rect 173791 94961 173839 94989
rect 173529 86175 173839 94961
rect 173529 86147 173577 86175
rect 173605 86147 173639 86175
rect 173667 86147 173701 86175
rect 173729 86147 173763 86175
rect 173791 86147 173839 86175
rect 173529 86113 173839 86147
rect 173529 86085 173577 86113
rect 173605 86085 173639 86113
rect 173667 86085 173701 86113
rect 173729 86085 173763 86113
rect 173791 86085 173839 86113
rect 173529 86051 173839 86085
rect 173529 86023 173577 86051
rect 173605 86023 173639 86051
rect 173667 86023 173701 86051
rect 173729 86023 173763 86051
rect 173791 86023 173839 86051
rect 173529 85989 173839 86023
rect 173529 85961 173577 85989
rect 173605 85961 173639 85989
rect 173667 85961 173701 85989
rect 173729 85961 173763 85989
rect 173791 85961 173839 85989
rect 173529 77175 173839 85961
rect 173529 77147 173577 77175
rect 173605 77147 173639 77175
rect 173667 77147 173701 77175
rect 173729 77147 173763 77175
rect 173791 77147 173839 77175
rect 173529 77113 173839 77147
rect 173529 77085 173577 77113
rect 173605 77085 173639 77113
rect 173667 77085 173701 77113
rect 173729 77085 173763 77113
rect 173791 77085 173839 77113
rect 173529 77051 173839 77085
rect 173529 77023 173577 77051
rect 173605 77023 173639 77051
rect 173667 77023 173701 77051
rect 173729 77023 173763 77051
rect 173791 77023 173839 77051
rect 173529 76989 173839 77023
rect 173529 76961 173577 76989
rect 173605 76961 173639 76989
rect 173667 76961 173701 76989
rect 173729 76961 173763 76989
rect 173791 76961 173839 76989
rect 173529 68175 173839 76961
rect 173529 68147 173577 68175
rect 173605 68147 173639 68175
rect 173667 68147 173701 68175
rect 173729 68147 173763 68175
rect 173791 68147 173839 68175
rect 173529 68113 173839 68147
rect 173529 68085 173577 68113
rect 173605 68085 173639 68113
rect 173667 68085 173701 68113
rect 173729 68085 173763 68113
rect 173791 68085 173839 68113
rect 173529 68051 173839 68085
rect 173529 68023 173577 68051
rect 173605 68023 173639 68051
rect 173667 68023 173701 68051
rect 173729 68023 173763 68051
rect 173791 68023 173839 68051
rect 173529 67989 173839 68023
rect 173529 67961 173577 67989
rect 173605 67961 173639 67989
rect 173667 67961 173701 67989
rect 173729 67961 173763 67989
rect 173791 67961 173839 67989
rect 173529 59175 173839 67961
rect 173529 59147 173577 59175
rect 173605 59147 173639 59175
rect 173667 59147 173701 59175
rect 173729 59147 173763 59175
rect 173791 59147 173839 59175
rect 173529 59113 173839 59147
rect 173529 59085 173577 59113
rect 173605 59085 173639 59113
rect 173667 59085 173701 59113
rect 173729 59085 173763 59113
rect 173791 59085 173839 59113
rect 173529 59051 173839 59085
rect 173529 59023 173577 59051
rect 173605 59023 173639 59051
rect 173667 59023 173701 59051
rect 173729 59023 173763 59051
rect 173791 59023 173839 59051
rect 173529 58989 173839 59023
rect 173529 58961 173577 58989
rect 173605 58961 173639 58989
rect 173667 58961 173701 58989
rect 173729 58961 173763 58989
rect 173791 58961 173839 58989
rect 173529 50175 173839 58961
rect 173529 50147 173577 50175
rect 173605 50147 173639 50175
rect 173667 50147 173701 50175
rect 173729 50147 173763 50175
rect 173791 50147 173839 50175
rect 173529 50113 173839 50147
rect 173529 50085 173577 50113
rect 173605 50085 173639 50113
rect 173667 50085 173701 50113
rect 173729 50085 173763 50113
rect 173791 50085 173839 50113
rect 173529 50051 173839 50085
rect 173529 50023 173577 50051
rect 173605 50023 173639 50051
rect 173667 50023 173701 50051
rect 173729 50023 173763 50051
rect 173791 50023 173839 50051
rect 173529 49989 173839 50023
rect 173529 49961 173577 49989
rect 173605 49961 173639 49989
rect 173667 49961 173701 49989
rect 173729 49961 173763 49989
rect 173791 49961 173839 49989
rect 173529 41175 173839 49961
rect 173529 41147 173577 41175
rect 173605 41147 173639 41175
rect 173667 41147 173701 41175
rect 173729 41147 173763 41175
rect 173791 41147 173839 41175
rect 173529 41113 173839 41147
rect 173529 41085 173577 41113
rect 173605 41085 173639 41113
rect 173667 41085 173701 41113
rect 173729 41085 173763 41113
rect 173791 41085 173839 41113
rect 173529 41051 173839 41085
rect 173529 41023 173577 41051
rect 173605 41023 173639 41051
rect 173667 41023 173701 41051
rect 173729 41023 173763 41051
rect 173791 41023 173839 41051
rect 173529 40989 173839 41023
rect 173529 40961 173577 40989
rect 173605 40961 173639 40989
rect 173667 40961 173701 40989
rect 173729 40961 173763 40989
rect 173791 40961 173839 40989
rect 173529 32175 173839 40961
rect 173529 32147 173577 32175
rect 173605 32147 173639 32175
rect 173667 32147 173701 32175
rect 173729 32147 173763 32175
rect 173791 32147 173839 32175
rect 173529 32113 173839 32147
rect 173529 32085 173577 32113
rect 173605 32085 173639 32113
rect 173667 32085 173701 32113
rect 173729 32085 173763 32113
rect 173791 32085 173839 32113
rect 173529 32051 173839 32085
rect 173529 32023 173577 32051
rect 173605 32023 173639 32051
rect 173667 32023 173701 32051
rect 173729 32023 173763 32051
rect 173791 32023 173839 32051
rect 173529 31989 173839 32023
rect 173529 31961 173577 31989
rect 173605 31961 173639 31989
rect 173667 31961 173701 31989
rect 173729 31961 173763 31989
rect 173791 31961 173839 31989
rect 173529 23175 173839 31961
rect 173529 23147 173577 23175
rect 173605 23147 173639 23175
rect 173667 23147 173701 23175
rect 173729 23147 173763 23175
rect 173791 23147 173839 23175
rect 173529 23113 173839 23147
rect 173529 23085 173577 23113
rect 173605 23085 173639 23113
rect 173667 23085 173701 23113
rect 173729 23085 173763 23113
rect 173791 23085 173839 23113
rect 173529 23051 173839 23085
rect 173529 23023 173577 23051
rect 173605 23023 173639 23051
rect 173667 23023 173701 23051
rect 173729 23023 173763 23051
rect 173791 23023 173839 23051
rect 173529 22989 173839 23023
rect 173529 22961 173577 22989
rect 173605 22961 173639 22989
rect 173667 22961 173701 22989
rect 173729 22961 173763 22989
rect 173791 22961 173839 22989
rect 173529 14175 173839 22961
rect 173529 14147 173577 14175
rect 173605 14147 173639 14175
rect 173667 14147 173701 14175
rect 173729 14147 173763 14175
rect 173791 14147 173839 14175
rect 173529 14113 173839 14147
rect 173529 14085 173577 14113
rect 173605 14085 173639 14113
rect 173667 14085 173701 14113
rect 173729 14085 173763 14113
rect 173791 14085 173839 14113
rect 173529 14051 173839 14085
rect 173529 14023 173577 14051
rect 173605 14023 173639 14051
rect 173667 14023 173701 14051
rect 173729 14023 173763 14051
rect 173791 14023 173839 14051
rect 173529 13989 173839 14023
rect 173529 13961 173577 13989
rect 173605 13961 173639 13989
rect 173667 13961 173701 13989
rect 173729 13961 173763 13989
rect 173791 13961 173839 13989
rect 173529 5175 173839 13961
rect 173529 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 173839 5175
rect 173529 5113 173839 5147
rect 173529 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 173839 5113
rect 173529 5051 173839 5085
rect 173529 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 173839 5051
rect 173529 4989 173839 5023
rect 173529 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 173839 4989
rect 173529 -560 173839 4961
rect 173529 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 173839 -560
rect 173529 -622 173839 -588
rect 173529 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 173839 -622
rect 173529 -684 173839 -650
rect 173529 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 173839 -684
rect 173529 -746 173839 -712
rect 173529 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 173839 -746
rect 173529 -822 173839 -774
rect 187029 92175 187339 100689
rect 187029 92147 187077 92175
rect 187105 92147 187139 92175
rect 187167 92147 187201 92175
rect 187229 92147 187263 92175
rect 187291 92147 187339 92175
rect 187029 92113 187339 92147
rect 187029 92085 187077 92113
rect 187105 92085 187139 92113
rect 187167 92085 187201 92113
rect 187229 92085 187263 92113
rect 187291 92085 187339 92113
rect 187029 92051 187339 92085
rect 187029 92023 187077 92051
rect 187105 92023 187139 92051
rect 187167 92023 187201 92051
rect 187229 92023 187263 92051
rect 187291 92023 187339 92051
rect 187029 91989 187339 92023
rect 187029 91961 187077 91989
rect 187105 91961 187139 91989
rect 187167 91961 187201 91989
rect 187229 91961 187263 91989
rect 187291 91961 187339 91989
rect 187029 83175 187339 91961
rect 187029 83147 187077 83175
rect 187105 83147 187139 83175
rect 187167 83147 187201 83175
rect 187229 83147 187263 83175
rect 187291 83147 187339 83175
rect 187029 83113 187339 83147
rect 187029 83085 187077 83113
rect 187105 83085 187139 83113
rect 187167 83085 187201 83113
rect 187229 83085 187263 83113
rect 187291 83085 187339 83113
rect 187029 83051 187339 83085
rect 187029 83023 187077 83051
rect 187105 83023 187139 83051
rect 187167 83023 187201 83051
rect 187229 83023 187263 83051
rect 187291 83023 187339 83051
rect 187029 82989 187339 83023
rect 187029 82961 187077 82989
rect 187105 82961 187139 82989
rect 187167 82961 187201 82989
rect 187229 82961 187263 82989
rect 187291 82961 187339 82989
rect 187029 74175 187339 82961
rect 187029 74147 187077 74175
rect 187105 74147 187139 74175
rect 187167 74147 187201 74175
rect 187229 74147 187263 74175
rect 187291 74147 187339 74175
rect 187029 74113 187339 74147
rect 187029 74085 187077 74113
rect 187105 74085 187139 74113
rect 187167 74085 187201 74113
rect 187229 74085 187263 74113
rect 187291 74085 187339 74113
rect 187029 74051 187339 74085
rect 187029 74023 187077 74051
rect 187105 74023 187139 74051
rect 187167 74023 187201 74051
rect 187229 74023 187263 74051
rect 187291 74023 187339 74051
rect 187029 73989 187339 74023
rect 187029 73961 187077 73989
rect 187105 73961 187139 73989
rect 187167 73961 187201 73989
rect 187229 73961 187263 73989
rect 187291 73961 187339 73989
rect 187029 65175 187339 73961
rect 187029 65147 187077 65175
rect 187105 65147 187139 65175
rect 187167 65147 187201 65175
rect 187229 65147 187263 65175
rect 187291 65147 187339 65175
rect 187029 65113 187339 65147
rect 187029 65085 187077 65113
rect 187105 65085 187139 65113
rect 187167 65085 187201 65113
rect 187229 65085 187263 65113
rect 187291 65085 187339 65113
rect 187029 65051 187339 65085
rect 187029 65023 187077 65051
rect 187105 65023 187139 65051
rect 187167 65023 187201 65051
rect 187229 65023 187263 65051
rect 187291 65023 187339 65051
rect 187029 64989 187339 65023
rect 187029 64961 187077 64989
rect 187105 64961 187139 64989
rect 187167 64961 187201 64989
rect 187229 64961 187263 64989
rect 187291 64961 187339 64989
rect 187029 56175 187339 64961
rect 187029 56147 187077 56175
rect 187105 56147 187139 56175
rect 187167 56147 187201 56175
rect 187229 56147 187263 56175
rect 187291 56147 187339 56175
rect 187029 56113 187339 56147
rect 187029 56085 187077 56113
rect 187105 56085 187139 56113
rect 187167 56085 187201 56113
rect 187229 56085 187263 56113
rect 187291 56085 187339 56113
rect 187029 56051 187339 56085
rect 187029 56023 187077 56051
rect 187105 56023 187139 56051
rect 187167 56023 187201 56051
rect 187229 56023 187263 56051
rect 187291 56023 187339 56051
rect 187029 55989 187339 56023
rect 187029 55961 187077 55989
rect 187105 55961 187139 55989
rect 187167 55961 187201 55989
rect 187229 55961 187263 55989
rect 187291 55961 187339 55989
rect 187029 47175 187339 55961
rect 187029 47147 187077 47175
rect 187105 47147 187139 47175
rect 187167 47147 187201 47175
rect 187229 47147 187263 47175
rect 187291 47147 187339 47175
rect 187029 47113 187339 47147
rect 187029 47085 187077 47113
rect 187105 47085 187139 47113
rect 187167 47085 187201 47113
rect 187229 47085 187263 47113
rect 187291 47085 187339 47113
rect 187029 47051 187339 47085
rect 187029 47023 187077 47051
rect 187105 47023 187139 47051
rect 187167 47023 187201 47051
rect 187229 47023 187263 47051
rect 187291 47023 187339 47051
rect 187029 46989 187339 47023
rect 187029 46961 187077 46989
rect 187105 46961 187139 46989
rect 187167 46961 187201 46989
rect 187229 46961 187263 46989
rect 187291 46961 187339 46989
rect 187029 38175 187339 46961
rect 187029 38147 187077 38175
rect 187105 38147 187139 38175
rect 187167 38147 187201 38175
rect 187229 38147 187263 38175
rect 187291 38147 187339 38175
rect 187029 38113 187339 38147
rect 187029 38085 187077 38113
rect 187105 38085 187139 38113
rect 187167 38085 187201 38113
rect 187229 38085 187263 38113
rect 187291 38085 187339 38113
rect 187029 38051 187339 38085
rect 187029 38023 187077 38051
rect 187105 38023 187139 38051
rect 187167 38023 187201 38051
rect 187229 38023 187263 38051
rect 187291 38023 187339 38051
rect 187029 37989 187339 38023
rect 187029 37961 187077 37989
rect 187105 37961 187139 37989
rect 187167 37961 187201 37989
rect 187229 37961 187263 37989
rect 187291 37961 187339 37989
rect 187029 29175 187339 37961
rect 187029 29147 187077 29175
rect 187105 29147 187139 29175
rect 187167 29147 187201 29175
rect 187229 29147 187263 29175
rect 187291 29147 187339 29175
rect 187029 29113 187339 29147
rect 187029 29085 187077 29113
rect 187105 29085 187139 29113
rect 187167 29085 187201 29113
rect 187229 29085 187263 29113
rect 187291 29085 187339 29113
rect 187029 29051 187339 29085
rect 187029 29023 187077 29051
rect 187105 29023 187139 29051
rect 187167 29023 187201 29051
rect 187229 29023 187263 29051
rect 187291 29023 187339 29051
rect 187029 28989 187339 29023
rect 187029 28961 187077 28989
rect 187105 28961 187139 28989
rect 187167 28961 187201 28989
rect 187229 28961 187263 28989
rect 187291 28961 187339 28989
rect 187029 20175 187339 28961
rect 187029 20147 187077 20175
rect 187105 20147 187139 20175
rect 187167 20147 187201 20175
rect 187229 20147 187263 20175
rect 187291 20147 187339 20175
rect 187029 20113 187339 20147
rect 187029 20085 187077 20113
rect 187105 20085 187139 20113
rect 187167 20085 187201 20113
rect 187229 20085 187263 20113
rect 187291 20085 187339 20113
rect 187029 20051 187339 20085
rect 187029 20023 187077 20051
rect 187105 20023 187139 20051
rect 187167 20023 187201 20051
rect 187229 20023 187263 20051
rect 187291 20023 187339 20051
rect 187029 19989 187339 20023
rect 187029 19961 187077 19989
rect 187105 19961 187139 19989
rect 187167 19961 187201 19989
rect 187229 19961 187263 19989
rect 187291 19961 187339 19989
rect 187029 11175 187339 19961
rect 187029 11147 187077 11175
rect 187105 11147 187139 11175
rect 187167 11147 187201 11175
rect 187229 11147 187263 11175
rect 187291 11147 187339 11175
rect 187029 11113 187339 11147
rect 187029 11085 187077 11113
rect 187105 11085 187139 11113
rect 187167 11085 187201 11113
rect 187229 11085 187263 11113
rect 187291 11085 187339 11113
rect 187029 11051 187339 11085
rect 187029 11023 187077 11051
rect 187105 11023 187139 11051
rect 187167 11023 187201 11051
rect 187229 11023 187263 11051
rect 187291 11023 187339 11051
rect 187029 10989 187339 11023
rect 187029 10961 187077 10989
rect 187105 10961 187139 10989
rect 187167 10961 187201 10989
rect 187229 10961 187263 10989
rect 187291 10961 187339 10989
rect 187029 2175 187339 10961
rect 187029 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 187339 2175
rect 187029 2113 187339 2147
rect 187029 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 187339 2113
rect 187029 2051 187339 2085
rect 187029 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 187339 2051
rect 187029 1989 187339 2023
rect 187029 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 187339 1989
rect 187029 -80 187339 1961
rect 187029 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 187339 -80
rect 187029 -142 187339 -108
rect 187029 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 187339 -142
rect 187029 -204 187339 -170
rect 187029 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 187339 -204
rect 187029 -266 187339 -232
rect 187029 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 187339 -266
rect 187029 -822 187339 -294
rect 188889 95175 189199 100689
rect 188889 95147 188937 95175
rect 188965 95147 188999 95175
rect 189027 95147 189061 95175
rect 189089 95147 189123 95175
rect 189151 95147 189199 95175
rect 188889 95113 189199 95147
rect 188889 95085 188937 95113
rect 188965 95085 188999 95113
rect 189027 95085 189061 95113
rect 189089 95085 189123 95113
rect 189151 95085 189199 95113
rect 188889 95051 189199 95085
rect 188889 95023 188937 95051
rect 188965 95023 188999 95051
rect 189027 95023 189061 95051
rect 189089 95023 189123 95051
rect 189151 95023 189199 95051
rect 188889 94989 189199 95023
rect 188889 94961 188937 94989
rect 188965 94961 188999 94989
rect 189027 94961 189061 94989
rect 189089 94961 189123 94989
rect 189151 94961 189199 94989
rect 188889 86175 189199 94961
rect 188889 86147 188937 86175
rect 188965 86147 188999 86175
rect 189027 86147 189061 86175
rect 189089 86147 189123 86175
rect 189151 86147 189199 86175
rect 188889 86113 189199 86147
rect 188889 86085 188937 86113
rect 188965 86085 188999 86113
rect 189027 86085 189061 86113
rect 189089 86085 189123 86113
rect 189151 86085 189199 86113
rect 188889 86051 189199 86085
rect 188889 86023 188937 86051
rect 188965 86023 188999 86051
rect 189027 86023 189061 86051
rect 189089 86023 189123 86051
rect 189151 86023 189199 86051
rect 188889 85989 189199 86023
rect 188889 85961 188937 85989
rect 188965 85961 188999 85989
rect 189027 85961 189061 85989
rect 189089 85961 189123 85989
rect 189151 85961 189199 85989
rect 188889 77175 189199 85961
rect 188889 77147 188937 77175
rect 188965 77147 188999 77175
rect 189027 77147 189061 77175
rect 189089 77147 189123 77175
rect 189151 77147 189199 77175
rect 188889 77113 189199 77147
rect 188889 77085 188937 77113
rect 188965 77085 188999 77113
rect 189027 77085 189061 77113
rect 189089 77085 189123 77113
rect 189151 77085 189199 77113
rect 188889 77051 189199 77085
rect 188889 77023 188937 77051
rect 188965 77023 188999 77051
rect 189027 77023 189061 77051
rect 189089 77023 189123 77051
rect 189151 77023 189199 77051
rect 188889 76989 189199 77023
rect 188889 76961 188937 76989
rect 188965 76961 188999 76989
rect 189027 76961 189061 76989
rect 189089 76961 189123 76989
rect 189151 76961 189199 76989
rect 188889 68175 189199 76961
rect 188889 68147 188937 68175
rect 188965 68147 188999 68175
rect 189027 68147 189061 68175
rect 189089 68147 189123 68175
rect 189151 68147 189199 68175
rect 188889 68113 189199 68147
rect 188889 68085 188937 68113
rect 188965 68085 188999 68113
rect 189027 68085 189061 68113
rect 189089 68085 189123 68113
rect 189151 68085 189199 68113
rect 188889 68051 189199 68085
rect 188889 68023 188937 68051
rect 188965 68023 188999 68051
rect 189027 68023 189061 68051
rect 189089 68023 189123 68051
rect 189151 68023 189199 68051
rect 188889 67989 189199 68023
rect 188889 67961 188937 67989
rect 188965 67961 188999 67989
rect 189027 67961 189061 67989
rect 189089 67961 189123 67989
rect 189151 67961 189199 67989
rect 188889 59175 189199 67961
rect 188889 59147 188937 59175
rect 188965 59147 188999 59175
rect 189027 59147 189061 59175
rect 189089 59147 189123 59175
rect 189151 59147 189199 59175
rect 188889 59113 189199 59147
rect 188889 59085 188937 59113
rect 188965 59085 188999 59113
rect 189027 59085 189061 59113
rect 189089 59085 189123 59113
rect 189151 59085 189199 59113
rect 188889 59051 189199 59085
rect 188889 59023 188937 59051
rect 188965 59023 188999 59051
rect 189027 59023 189061 59051
rect 189089 59023 189123 59051
rect 189151 59023 189199 59051
rect 188889 58989 189199 59023
rect 188889 58961 188937 58989
rect 188965 58961 188999 58989
rect 189027 58961 189061 58989
rect 189089 58961 189123 58989
rect 189151 58961 189199 58989
rect 188889 50175 189199 58961
rect 188889 50147 188937 50175
rect 188965 50147 188999 50175
rect 189027 50147 189061 50175
rect 189089 50147 189123 50175
rect 189151 50147 189199 50175
rect 188889 50113 189199 50147
rect 188889 50085 188937 50113
rect 188965 50085 188999 50113
rect 189027 50085 189061 50113
rect 189089 50085 189123 50113
rect 189151 50085 189199 50113
rect 188889 50051 189199 50085
rect 188889 50023 188937 50051
rect 188965 50023 188999 50051
rect 189027 50023 189061 50051
rect 189089 50023 189123 50051
rect 189151 50023 189199 50051
rect 188889 49989 189199 50023
rect 188889 49961 188937 49989
rect 188965 49961 188999 49989
rect 189027 49961 189061 49989
rect 189089 49961 189123 49989
rect 189151 49961 189199 49989
rect 188889 41175 189199 49961
rect 188889 41147 188937 41175
rect 188965 41147 188999 41175
rect 189027 41147 189061 41175
rect 189089 41147 189123 41175
rect 189151 41147 189199 41175
rect 188889 41113 189199 41147
rect 188889 41085 188937 41113
rect 188965 41085 188999 41113
rect 189027 41085 189061 41113
rect 189089 41085 189123 41113
rect 189151 41085 189199 41113
rect 188889 41051 189199 41085
rect 188889 41023 188937 41051
rect 188965 41023 188999 41051
rect 189027 41023 189061 41051
rect 189089 41023 189123 41051
rect 189151 41023 189199 41051
rect 188889 40989 189199 41023
rect 188889 40961 188937 40989
rect 188965 40961 188999 40989
rect 189027 40961 189061 40989
rect 189089 40961 189123 40989
rect 189151 40961 189199 40989
rect 188889 32175 189199 40961
rect 188889 32147 188937 32175
rect 188965 32147 188999 32175
rect 189027 32147 189061 32175
rect 189089 32147 189123 32175
rect 189151 32147 189199 32175
rect 188889 32113 189199 32147
rect 188889 32085 188937 32113
rect 188965 32085 188999 32113
rect 189027 32085 189061 32113
rect 189089 32085 189123 32113
rect 189151 32085 189199 32113
rect 188889 32051 189199 32085
rect 188889 32023 188937 32051
rect 188965 32023 188999 32051
rect 189027 32023 189061 32051
rect 189089 32023 189123 32051
rect 189151 32023 189199 32051
rect 188889 31989 189199 32023
rect 188889 31961 188937 31989
rect 188965 31961 188999 31989
rect 189027 31961 189061 31989
rect 189089 31961 189123 31989
rect 189151 31961 189199 31989
rect 188889 23175 189199 31961
rect 188889 23147 188937 23175
rect 188965 23147 188999 23175
rect 189027 23147 189061 23175
rect 189089 23147 189123 23175
rect 189151 23147 189199 23175
rect 188889 23113 189199 23147
rect 188889 23085 188937 23113
rect 188965 23085 188999 23113
rect 189027 23085 189061 23113
rect 189089 23085 189123 23113
rect 189151 23085 189199 23113
rect 188889 23051 189199 23085
rect 188889 23023 188937 23051
rect 188965 23023 188999 23051
rect 189027 23023 189061 23051
rect 189089 23023 189123 23051
rect 189151 23023 189199 23051
rect 188889 22989 189199 23023
rect 188889 22961 188937 22989
rect 188965 22961 188999 22989
rect 189027 22961 189061 22989
rect 189089 22961 189123 22989
rect 189151 22961 189199 22989
rect 188889 14175 189199 22961
rect 188889 14147 188937 14175
rect 188965 14147 188999 14175
rect 189027 14147 189061 14175
rect 189089 14147 189123 14175
rect 189151 14147 189199 14175
rect 188889 14113 189199 14147
rect 188889 14085 188937 14113
rect 188965 14085 188999 14113
rect 189027 14085 189061 14113
rect 189089 14085 189123 14113
rect 189151 14085 189199 14113
rect 188889 14051 189199 14085
rect 188889 14023 188937 14051
rect 188965 14023 188999 14051
rect 189027 14023 189061 14051
rect 189089 14023 189123 14051
rect 189151 14023 189199 14051
rect 188889 13989 189199 14023
rect 188889 13961 188937 13989
rect 188965 13961 188999 13989
rect 189027 13961 189061 13989
rect 189089 13961 189123 13989
rect 189151 13961 189199 13989
rect 188889 5175 189199 13961
rect 188889 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 189199 5175
rect 188889 5113 189199 5147
rect 188889 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 189199 5113
rect 188889 5051 189199 5085
rect 188889 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 189199 5051
rect 188889 4989 189199 5023
rect 188889 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 189199 4989
rect 188889 -560 189199 4961
rect 188889 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 189199 -560
rect 188889 -622 189199 -588
rect 188889 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 189199 -622
rect 188889 -684 189199 -650
rect 188889 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 189199 -684
rect 188889 -746 189199 -712
rect 188889 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 189199 -746
rect 188889 -822 189199 -774
rect 202389 92175 202699 100689
rect 202389 92147 202437 92175
rect 202465 92147 202499 92175
rect 202527 92147 202561 92175
rect 202589 92147 202623 92175
rect 202651 92147 202699 92175
rect 202389 92113 202699 92147
rect 202389 92085 202437 92113
rect 202465 92085 202499 92113
rect 202527 92085 202561 92113
rect 202589 92085 202623 92113
rect 202651 92085 202699 92113
rect 202389 92051 202699 92085
rect 202389 92023 202437 92051
rect 202465 92023 202499 92051
rect 202527 92023 202561 92051
rect 202589 92023 202623 92051
rect 202651 92023 202699 92051
rect 202389 91989 202699 92023
rect 202389 91961 202437 91989
rect 202465 91961 202499 91989
rect 202527 91961 202561 91989
rect 202589 91961 202623 91989
rect 202651 91961 202699 91989
rect 202389 83175 202699 91961
rect 202389 83147 202437 83175
rect 202465 83147 202499 83175
rect 202527 83147 202561 83175
rect 202589 83147 202623 83175
rect 202651 83147 202699 83175
rect 202389 83113 202699 83147
rect 202389 83085 202437 83113
rect 202465 83085 202499 83113
rect 202527 83085 202561 83113
rect 202589 83085 202623 83113
rect 202651 83085 202699 83113
rect 202389 83051 202699 83085
rect 202389 83023 202437 83051
rect 202465 83023 202499 83051
rect 202527 83023 202561 83051
rect 202589 83023 202623 83051
rect 202651 83023 202699 83051
rect 202389 82989 202699 83023
rect 202389 82961 202437 82989
rect 202465 82961 202499 82989
rect 202527 82961 202561 82989
rect 202589 82961 202623 82989
rect 202651 82961 202699 82989
rect 202389 74175 202699 82961
rect 202389 74147 202437 74175
rect 202465 74147 202499 74175
rect 202527 74147 202561 74175
rect 202589 74147 202623 74175
rect 202651 74147 202699 74175
rect 202389 74113 202699 74147
rect 202389 74085 202437 74113
rect 202465 74085 202499 74113
rect 202527 74085 202561 74113
rect 202589 74085 202623 74113
rect 202651 74085 202699 74113
rect 202389 74051 202699 74085
rect 202389 74023 202437 74051
rect 202465 74023 202499 74051
rect 202527 74023 202561 74051
rect 202589 74023 202623 74051
rect 202651 74023 202699 74051
rect 202389 73989 202699 74023
rect 202389 73961 202437 73989
rect 202465 73961 202499 73989
rect 202527 73961 202561 73989
rect 202589 73961 202623 73989
rect 202651 73961 202699 73989
rect 202389 65175 202699 73961
rect 202389 65147 202437 65175
rect 202465 65147 202499 65175
rect 202527 65147 202561 65175
rect 202589 65147 202623 65175
rect 202651 65147 202699 65175
rect 202389 65113 202699 65147
rect 202389 65085 202437 65113
rect 202465 65085 202499 65113
rect 202527 65085 202561 65113
rect 202589 65085 202623 65113
rect 202651 65085 202699 65113
rect 202389 65051 202699 65085
rect 202389 65023 202437 65051
rect 202465 65023 202499 65051
rect 202527 65023 202561 65051
rect 202589 65023 202623 65051
rect 202651 65023 202699 65051
rect 202389 64989 202699 65023
rect 202389 64961 202437 64989
rect 202465 64961 202499 64989
rect 202527 64961 202561 64989
rect 202589 64961 202623 64989
rect 202651 64961 202699 64989
rect 202389 56175 202699 64961
rect 202389 56147 202437 56175
rect 202465 56147 202499 56175
rect 202527 56147 202561 56175
rect 202589 56147 202623 56175
rect 202651 56147 202699 56175
rect 202389 56113 202699 56147
rect 202389 56085 202437 56113
rect 202465 56085 202499 56113
rect 202527 56085 202561 56113
rect 202589 56085 202623 56113
rect 202651 56085 202699 56113
rect 202389 56051 202699 56085
rect 202389 56023 202437 56051
rect 202465 56023 202499 56051
rect 202527 56023 202561 56051
rect 202589 56023 202623 56051
rect 202651 56023 202699 56051
rect 202389 55989 202699 56023
rect 202389 55961 202437 55989
rect 202465 55961 202499 55989
rect 202527 55961 202561 55989
rect 202589 55961 202623 55989
rect 202651 55961 202699 55989
rect 202389 47175 202699 55961
rect 202389 47147 202437 47175
rect 202465 47147 202499 47175
rect 202527 47147 202561 47175
rect 202589 47147 202623 47175
rect 202651 47147 202699 47175
rect 202389 47113 202699 47147
rect 202389 47085 202437 47113
rect 202465 47085 202499 47113
rect 202527 47085 202561 47113
rect 202589 47085 202623 47113
rect 202651 47085 202699 47113
rect 202389 47051 202699 47085
rect 202389 47023 202437 47051
rect 202465 47023 202499 47051
rect 202527 47023 202561 47051
rect 202589 47023 202623 47051
rect 202651 47023 202699 47051
rect 202389 46989 202699 47023
rect 202389 46961 202437 46989
rect 202465 46961 202499 46989
rect 202527 46961 202561 46989
rect 202589 46961 202623 46989
rect 202651 46961 202699 46989
rect 202389 38175 202699 46961
rect 202389 38147 202437 38175
rect 202465 38147 202499 38175
rect 202527 38147 202561 38175
rect 202589 38147 202623 38175
rect 202651 38147 202699 38175
rect 202389 38113 202699 38147
rect 202389 38085 202437 38113
rect 202465 38085 202499 38113
rect 202527 38085 202561 38113
rect 202589 38085 202623 38113
rect 202651 38085 202699 38113
rect 202389 38051 202699 38085
rect 202389 38023 202437 38051
rect 202465 38023 202499 38051
rect 202527 38023 202561 38051
rect 202589 38023 202623 38051
rect 202651 38023 202699 38051
rect 202389 37989 202699 38023
rect 202389 37961 202437 37989
rect 202465 37961 202499 37989
rect 202527 37961 202561 37989
rect 202589 37961 202623 37989
rect 202651 37961 202699 37989
rect 202389 29175 202699 37961
rect 202389 29147 202437 29175
rect 202465 29147 202499 29175
rect 202527 29147 202561 29175
rect 202589 29147 202623 29175
rect 202651 29147 202699 29175
rect 202389 29113 202699 29147
rect 202389 29085 202437 29113
rect 202465 29085 202499 29113
rect 202527 29085 202561 29113
rect 202589 29085 202623 29113
rect 202651 29085 202699 29113
rect 202389 29051 202699 29085
rect 202389 29023 202437 29051
rect 202465 29023 202499 29051
rect 202527 29023 202561 29051
rect 202589 29023 202623 29051
rect 202651 29023 202699 29051
rect 202389 28989 202699 29023
rect 202389 28961 202437 28989
rect 202465 28961 202499 28989
rect 202527 28961 202561 28989
rect 202589 28961 202623 28989
rect 202651 28961 202699 28989
rect 202389 20175 202699 28961
rect 202389 20147 202437 20175
rect 202465 20147 202499 20175
rect 202527 20147 202561 20175
rect 202589 20147 202623 20175
rect 202651 20147 202699 20175
rect 202389 20113 202699 20147
rect 202389 20085 202437 20113
rect 202465 20085 202499 20113
rect 202527 20085 202561 20113
rect 202589 20085 202623 20113
rect 202651 20085 202699 20113
rect 202389 20051 202699 20085
rect 202389 20023 202437 20051
rect 202465 20023 202499 20051
rect 202527 20023 202561 20051
rect 202589 20023 202623 20051
rect 202651 20023 202699 20051
rect 202389 19989 202699 20023
rect 202389 19961 202437 19989
rect 202465 19961 202499 19989
rect 202527 19961 202561 19989
rect 202589 19961 202623 19989
rect 202651 19961 202699 19989
rect 202389 11175 202699 19961
rect 202389 11147 202437 11175
rect 202465 11147 202499 11175
rect 202527 11147 202561 11175
rect 202589 11147 202623 11175
rect 202651 11147 202699 11175
rect 202389 11113 202699 11147
rect 202389 11085 202437 11113
rect 202465 11085 202499 11113
rect 202527 11085 202561 11113
rect 202589 11085 202623 11113
rect 202651 11085 202699 11113
rect 202389 11051 202699 11085
rect 202389 11023 202437 11051
rect 202465 11023 202499 11051
rect 202527 11023 202561 11051
rect 202589 11023 202623 11051
rect 202651 11023 202699 11051
rect 202389 10989 202699 11023
rect 202389 10961 202437 10989
rect 202465 10961 202499 10989
rect 202527 10961 202561 10989
rect 202589 10961 202623 10989
rect 202651 10961 202699 10989
rect 202389 2175 202699 10961
rect 202389 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 202699 2175
rect 202389 2113 202699 2147
rect 202389 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 202699 2113
rect 202389 2051 202699 2085
rect 202389 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 202699 2051
rect 202389 1989 202699 2023
rect 202389 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 202699 1989
rect 202389 -80 202699 1961
rect 202389 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 202699 -80
rect 202389 -142 202699 -108
rect 202389 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 202699 -142
rect 202389 -204 202699 -170
rect 202389 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 202699 -204
rect 202389 -266 202699 -232
rect 202389 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 202699 -266
rect 202389 -822 202699 -294
rect 204249 95175 204559 100689
rect 204249 95147 204297 95175
rect 204325 95147 204359 95175
rect 204387 95147 204421 95175
rect 204449 95147 204483 95175
rect 204511 95147 204559 95175
rect 204249 95113 204559 95147
rect 204249 95085 204297 95113
rect 204325 95085 204359 95113
rect 204387 95085 204421 95113
rect 204449 95085 204483 95113
rect 204511 95085 204559 95113
rect 204249 95051 204559 95085
rect 204249 95023 204297 95051
rect 204325 95023 204359 95051
rect 204387 95023 204421 95051
rect 204449 95023 204483 95051
rect 204511 95023 204559 95051
rect 204249 94989 204559 95023
rect 204249 94961 204297 94989
rect 204325 94961 204359 94989
rect 204387 94961 204421 94989
rect 204449 94961 204483 94989
rect 204511 94961 204559 94989
rect 204249 86175 204559 94961
rect 204249 86147 204297 86175
rect 204325 86147 204359 86175
rect 204387 86147 204421 86175
rect 204449 86147 204483 86175
rect 204511 86147 204559 86175
rect 204249 86113 204559 86147
rect 204249 86085 204297 86113
rect 204325 86085 204359 86113
rect 204387 86085 204421 86113
rect 204449 86085 204483 86113
rect 204511 86085 204559 86113
rect 204249 86051 204559 86085
rect 204249 86023 204297 86051
rect 204325 86023 204359 86051
rect 204387 86023 204421 86051
rect 204449 86023 204483 86051
rect 204511 86023 204559 86051
rect 204249 85989 204559 86023
rect 204249 85961 204297 85989
rect 204325 85961 204359 85989
rect 204387 85961 204421 85989
rect 204449 85961 204483 85989
rect 204511 85961 204559 85989
rect 204249 77175 204559 85961
rect 204249 77147 204297 77175
rect 204325 77147 204359 77175
rect 204387 77147 204421 77175
rect 204449 77147 204483 77175
rect 204511 77147 204559 77175
rect 204249 77113 204559 77147
rect 204249 77085 204297 77113
rect 204325 77085 204359 77113
rect 204387 77085 204421 77113
rect 204449 77085 204483 77113
rect 204511 77085 204559 77113
rect 204249 77051 204559 77085
rect 204249 77023 204297 77051
rect 204325 77023 204359 77051
rect 204387 77023 204421 77051
rect 204449 77023 204483 77051
rect 204511 77023 204559 77051
rect 204249 76989 204559 77023
rect 204249 76961 204297 76989
rect 204325 76961 204359 76989
rect 204387 76961 204421 76989
rect 204449 76961 204483 76989
rect 204511 76961 204559 76989
rect 204249 68175 204559 76961
rect 204249 68147 204297 68175
rect 204325 68147 204359 68175
rect 204387 68147 204421 68175
rect 204449 68147 204483 68175
rect 204511 68147 204559 68175
rect 204249 68113 204559 68147
rect 204249 68085 204297 68113
rect 204325 68085 204359 68113
rect 204387 68085 204421 68113
rect 204449 68085 204483 68113
rect 204511 68085 204559 68113
rect 204249 68051 204559 68085
rect 204249 68023 204297 68051
rect 204325 68023 204359 68051
rect 204387 68023 204421 68051
rect 204449 68023 204483 68051
rect 204511 68023 204559 68051
rect 204249 67989 204559 68023
rect 204249 67961 204297 67989
rect 204325 67961 204359 67989
rect 204387 67961 204421 67989
rect 204449 67961 204483 67989
rect 204511 67961 204559 67989
rect 204249 59175 204559 67961
rect 204249 59147 204297 59175
rect 204325 59147 204359 59175
rect 204387 59147 204421 59175
rect 204449 59147 204483 59175
rect 204511 59147 204559 59175
rect 204249 59113 204559 59147
rect 204249 59085 204297 59113
rect 204325 59085 204359 59113
rect 204387 59085 204421 59113
rect 204449 59085 204483 59113
rect 204511 59085 204559 59113
rect 204249 59051 204559 59085
rect 204249 59023 204297 59051
rect 204325 59023 204359 59051
rect 204387 59023 204421 59051
rect 204449 59023 204483 59051
rect 204511 59023 204559 59051
rect 204249 58989 204559 59023
rect 204249 58961 204297 58989
rect 204325 58961 204359 58989
rect 204387 58961 204421 58989
rect 204449 58961 204483 58989
rect 204511 58961 204559 58989
rect 204249 50175 204559 58961
rect 204249 50147 204297 50175
rect 204325 50147 204359 50175
rect 204387 50147 204421 50175
rect 204449 50147 204483 50175
rect 204511 50147 204559 50175
rect 204249 50113 204559 50147
rect 204249 50085 204297 50113
rect 204325 50085 204359 50113
rect 204387 50085 204421 50113
rect 204449 50085 204483 50113
rect 204511 50085 204559 50113
rect 204249 50051 204559 50085
rect 204249 50023 204297 50051
rect 204325 50023 204359 50051
rect 204387 50023 204421 50051
rect 204449 50023 204483 50051
rect 204511 50023 204559 50051
rect 204249 49989 204559 50023
rect 204249 49961 204297 49989
rect 204325 49961 204359 49989
rect 204387 49961 204421 49989
rect 204449 49961 204483 49989
rect 204511 49961 204559 49989
rect 204249 41175 204559 49961
rect 204249 41147 204297 41175
rect 204325 41147 204359 41175
rect 204387 41147 204421 41175
rect 204449 41147 204483 41175
rect 204511 41147 204559 41175
rect 204249 41113 204559 41147
rect 204249 41085 204297 41113
rect 204325 41085 204359 41113
rect 204387 41085 204421 41113
rect 204449 41085 204483 41113
rect 204511 41085 204559 41113
rect 204249 41051 204559 41085
rect 204249 41023 204297 41051
rect 204325 41023 204359 41051
rect 204387 41023 204421 41051
rect 204449 41023 204483 41051
rect 204511 41023 204559 41051
rect 204249 40989 204559 41023
rect 204249 40961 204297 40989
rect 204325 40961 204359 40989
rect 204387 40961 204421 40989
rect 204449 40961 204483 40989
rect 204511 40961 204559 40989
rect 204249 32175 204559 40961
rect 204249 32147 204297 32175
rect 204325 32147 204359 32175
rect 204387 32147 204421 32175
rect 204449 32147 204483 32175
rect 204511 32147 204559 32175
rect 204249 32113 204559 32147
rect 204249 32085 204297 32113
rect 204325 32085 204359 32113
rect 204387 32085 204421 32113
rect 204449 32085 204483 32113
rect 204511 32085 204559 32113
rect 204249 32051 204559 32085
rect 204249 32023 204297 32051
rect 204325 32023 204359 32051
rect 204387 32023 204421 32051
rect 204449 32023 204483 32051
rect 204511 32023 204559 32051
rect 204249 31989 204559 32023
rect 204249 31961 204297 31989
rect 204325 31961 204359 31989
rect 204387 31961 204421 31989
rect 204449 31961 204483 31989
rect 204511 31961 204559 31989
rect 204249 23175 204559 31961
rect 204249 23147 204297 23175
rect 204325 23147 204359 23175
rect 204387 23147 204421 23175
rect 204449 23147 204483 23175
rect 204511 23147 204559 23175
rect 204249 23113 204559 23147
rect 204249 23085 204297 23113
rect 204325 23085 204359 23113
rect 204387 23085 204421 23113
rect 204449 23085 204483 23113
rect 204511 23085 204559 23113
rect 204249 23051 204559 23085
rect 204249 23023 204297 23051
rect 204325 23023 204359 23051
rect 204387 23023 204421 23051
rect 204449 23023 204483 23051
rect 204511 23023 204559 23051
rect 204249 22989 204559 23023
rect 204249 22961 204297 22989
rect 204325 22961 204359 22989
rect 204387 22961 204421 22989
rect 204449 22961 204483 22989
rect 204511 22961 204559 22989
rect 204249 14175 204559 22961
rect 204249 14147 204297 14175
rect 204325 14147 204359 14175
rect 204387 14147 204421 14175
rect 204449 14147 204483 14175
rect 204511 14147 204559 14175
rect 204249 14113 204559 14147
rect 204249 14085 204297 14113
rect 204325 14085 204359 14113
rect 204387 14085 204421 14113
rect 204449 14085 204483 14113
rect 204511 14085 204559 14113
rect 204249 14051 204559 14085
rect 204249 14023 204297 14051
rect 204325 14023 204359 14051
rect 204387 14023 204421 14051
rect 204449 14023 204483 14051
rect 204511 14023 204559 14051
rect 204249 13989 204559 14023
rect 204249 13961 204297 13989
rect 204325 13961 204359 13989
rect 204387 13961 204421 13989
rect 204449 13961 204483 13989
rect 204511 13961 204559 13989
rect 204249 5175 204559 13961
rect 204249 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 204559 5175
rect 204249 5113 204559 5147
rect 204249 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 204559 5113
rect 204249 5051 204559 5085
rect 204249 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 204559 5051
rect 204249 4989 204559 5023
rect 204249 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 204559 4989
rect 204249 -560 204559 4961
rect 204249 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 204559 -560
rect 204249 -622 204559 -588
rect 204249 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 204559 -622
rect 204249 -684 204559 -650
rect 204249 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 204559 -684
rect 204249 -746 204559 -712
rect 204249 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 204559 -746
rect 204249 -822 204559 -774
rect 217749 92175 218059 100689
rect 217749 92147 217797 92175
rect 217825 92147 217859 92175
rect 217887 92147 217921 92175
rect 217949 92147 217983 92175
rect 218011 92147 218059 92175
rect 217749 92113 218059 92147
rect 217749 92085 217797 92113
rect 217825 92085 217859 92113
rect 217887 92085 217921 92113
rect 217949 92085 217983 92113
rect 218011 92085 218059 92113
rect 217749 92051 218059 92085
rect 217749 92023 217797 92051
rect 217825 92023 217859 92051
rect 217887 92023 217921 92051
rect 217949 92023 217983 92051
rect 218011 92023 218059 92051
rect 217749 91989 218059 92023
rect 217749 91961 217797 91989
rect 217825 91961 217859 91989
rect 217887 91961 217921 91989
rect 217949 91961 217983 91989
rect 218011 91961 218059 91989
rect 217749 83175 218059 91961
rect 217749 83147 217797 83175
rect 217825 83147 217859 83175
rect 217887 83147 217921 83175
rect 217949 83147 217983 83175
rect 218011 83147 218059 83175
rect 217749 83113 218059 83147
rect 217749 83085 217797 83113
rect 217825 83085 217859 83113
rect 217887 83085 217921 83113
rect 217949 83085 217983 83113
rect 218011 83085 218059 83113
rect 217749 83051 218059 83085
rect 217749 83023 217797 83051
rect 217825 83023 217859 83051
rect 217887 83023 217921 83051
rect 217949 83023 217983 83051
rect 218011 83023 218059 83051
rect 217749 82989 218059 83023
rect 217749 82961 217797 82989
rect 217825 82961 217859 82989
rect 217887 82961 217921 82989
rect 217949 82961 217983 82989
rect 218011 82961 218059 82989
rect 217749 74175 218059 82961
rect 217749 74147 217797 74175
rect 217825 74147 217859 74175
rect 217887 74147 217921 74175
rect 217949 74147 217983 74175
rect 218011 74147 218059 74175
rect 217749 74113 218059 74147
rect 217749 74085 217797 74113
rect 217825 74085 217859 74113
rect 217887 74085 217921 74113
rect 217949 74085 217983 74113
rect 218011 74085 218059 74113
rect 217749 74051 218059 74085
rect 217749 74023 217797 74051
rect 217825 74023 217859 74051
rect 217887 74023 217921 74051
rect 217949 74023 217983 74051
rect 218011 74023 218059 74051
rect 217749 73989 218059 74023
rect 217749 73961 217797 73989
rect 217825 73961 217859 73989
rect 217887 73961 217921 73989
rect 217949 73961 217983 73989
rect 218011 73961 218059 73989
rect 217749 65175 218059 73961
rect 217749 65147 217797 65175
rect 217825 65147 217859 65175
rect 217887 65147 217921 65175
rect 217949 65147 217983 65175
rect 218011 65147 218059 65175
rect 217749 65113 218059 65147
rect 217749 65085 217797 65113
rect 217825 65085 217859 65113
rect 217887 65085 217921 65113
rect 217949 65085 217983 65113
rect 218011 65085 218059 65113
rect 217749 65051 218059 65085
rect 217749 65023 217797 65051
rect 217825 65023 217859 65051
rect 217887 65023 217921 65051
rect 217949 65023 217983 65051
rect 218011 65023 218059 65051
rect 217749 64989 218059 65023
rect 217749 64961 217797 64989
rect 217825 64961 217859 64989
rect 217887 64961 217921 64989
rect 217949 64961 217983 64989
rect 218011 64961 218059 64989
rect 217749 56175 218059 64961
rect 217749 56147 217797 56175
rect 217825 56147 217859 56175
rect 217887 56147 217921 56175
rect 217949 56147 217983 56175
rect 218011 56147 218059 56175
rect 217749 56113 218059 56147
rect 217749 56085 217797 56113
rect 217825 56085 217859 56113
rect 217887 56085 217921 56113
rect 217949 56085 217983 56113
rect 218011 56085 218059 56113
rect 217749 56051 218059 56085
rect 217749 56023 217797 56051
rect 217825 56023 217859 56051
rect 217887 56023 217921 56051
rect 217949 56023 217983 56051
rect 218011 56023 218059 56051
rect 217749 55989 218059 56023
rect 217749 55961 217797 55989
rect 217825 55961 217859 55989
rect 217887 55961 217921 55989
rect 217949 55961 217983 55989
rect 218011 55961 218059 55989
rect 217749 47175 218059 55961
rect 217749 47147 217797 47175
rect 217825 47147 217859 47175
rect 217887 47147 217921 47175
rect 217949 47147 217983 47175
rect 218011 47147 218059 47175
rect 217749 47113 218059 47147
rect 217749 47085 217797 47113
rect 217825 47085 217859 47113
rect 217887 47085 217921 47113
rect 217949 47085 217983 47113
rect 218011 47085 218059 47113
rect 217749 47051 218059 47085
rect 217749 47023 217797 47051
rect 217825 47023 217859 47051
rect 217887 47023 217921 47051
rect 217949 47023 217983 47051
rect 218011 47023 218059 47051
rect 217749 46989 218059 47023
rect 217749 46961 217797 46989
rect 217825 46961 217859 46989
rect 217887 46961 217921 46989
rect 217949 46961 217983 46989
rect 218011 46961 218059 46989
rect 217749 38175 218059 46961
rect 217749 38147 217797 38175
rect 217825 38147 217859 38175
rect 217887 38147 217921 38175
rect 217949 38147 217983 38175
rect 218011 38147 218059 38175
rect 217749 38113 218059 38147
rect 217749 38085 217797 38113
rect 217825 38085 217859 38113
rect 217887 38085 217921 38113
rect 217949 38085 217983 38113
rect 218011 38085 218059 38113
rect 217749 38051 218059 38085
rect 217749 38023 217797 38051
rect 217825 38023 217859 38051
rect 217887 38023 217921 38051
rect 217949 38023 217983 38051
rect 218011 38023 218059 38051
rect 217749 37989 218059 38023
rect 217749 37961 217797 37989
rect 217825 37961 217859 37989
rect 217887 37961 217921 37989
rect 217949 37961 217983 37989
rect 218011 37961 218059 37989
rect 217749 29175 218059 37961
rect 217749 29147 217797 29175
rect 217825 29147 217859 29175
rect 217887 29147 217921 29175
rect 217949 29147 217983 29175
rect 218011 29147 218059 29175
rect 217749 29113 218059 29147
rect 217749 29085 217797 29113
rect 217825 29085 217859 29113
rect 217887 29085 217921 29113
rect 217949 29085 217983 29113
rect 218011 29085 218059 29113
rect 217749 29051 218059 29085
rect 217749 29023 217797 29051
rect 217825 29023 217859 29051
rect 217887 29023 217921 29051
rect 217949 29023 217983 29051
rect 218011 29023 218059 29051
rect 217749 28989 218059 29023
rect 217749 28961 217797 28989
rect 217825 28961 217859 28989
rect 217887 28961 217921 28989
rect 217949 28961 217983 28989
rect 218011 28961 218059 28989
rect 217749 20175 218059 28961
rect 217749 20147 217797 20175
rect 217825 20147 217859 20175
rect 217887 20147 217921 20175
rect 217949 20147 217983 20175
rect 218011 20147 218059 20175
rect 217749 20113 218059 20147
rect 217749 20085 217797 20113
rect 217825 20085 217859 20113
rect 217887 20085 217921 20113
rect 217949 20085 217983 20113
rect 218011 20085 218059 20113
rect 217749 20051 218059 20085
rect 217749 20023 217797 20051
rect 217825 20023 217859 20051
rect 217887 20023 217921 20051
rect 217949 20023 217983 20051
rect 218011 20023 218059 20051
rect 217749 19989 218059 20023
rect 217749 19961 217797 19989
rect 217825 19961 217859 19989
rect 217887 19961 217921 19989
rect 217949 19961 217983 19989
rect 218011 19961 218059 19989
rect 217749 11175 218059 19961
rect 217749 11147 217797 11175
rect 217825 11147 217859 11175
rect 217887 11147 217921 11175
rect 217949 11147 217983 11175
rect 218011 11147 218059 11175
rect 217749 11113 218059 11147
rect 217749 11085 217797 11113
rect 217825 11085 217859 11113
rect 217887 11085 217921 11113
rect 217949 11085 217983 11113
rect 218011 11085 218059 11113
rect 217749 11051 218059 11085
rect 217749 11023 217797 11051
rect 217825 11023 217859 11051
rect 217887 11023 217921 11051
rect 217949 11023 217983 11051
rect 218011 11023 218059 11051
rect 217749 10989 218059 11023
rect 217749 10961 217797 10989
rect 217825 10961 217859 10989
rect 217887 10961 217921 10989
rect 217949 10961 217983 10989
rect 218011 10961 218059 10989
rect 217749 2175 218059 10961
rect 217749 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 218059 2175
rect 217749 2113 218059 2147
rect 217749 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 218059 2113
rect 217749 2051 218059 2085
rect 217749 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 218059 2051
rect 217749 1989 218059 2023
rect 217749 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 218059 1989
rect 217749 -80 218059 1961
rect 217749 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 218059 -80
rect 217749 -142 218059 -108
rect 217749 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 218059 -142
rect 217749 -204 218059 -170
rect 217749 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 218059 -204
rect 217749 -266 218059 -232
rect 217749 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 218059 -266
rect 217749 -822 218059 -294
rect 219609 95175 219919 100689
rect 219609 95147 219657 95175
rect 219685 95147 219719 95175
rect 219747 95147 219781 95175
rect 219809 95147 219843 95175
rect 219871 95147 219919 95175
rect 219609 95113 219919 95147
rect 219609 95085 219657 95113
rect 219685 95085 219719 95113
rect 219747 95085 219781 95113
rect 219809 95085 219843 95113
rect 219871 95085 219919 95113
rect 219609 95051 219919 95085
rect 219609 95023 219657 95051
rect 219685 95023 219719 95051
rect 219747 95023 219781 95051
rect 219809 95023 219843 95051
rect 219871 95023 219919 95051
rect 219609 94989 219919 95023
rect 219609 94961 219657 94989
rect 219685 94961 219719 94989
rect 219747 94961 219781 94989
rect 219809 94961 219843 94989
rect 219871 94961 219919 94989
rect 219609 86175 219919 94961
rect 219609 86147 219657 86175
rect 219685 86147 219719 86175
rect 219747 86147 219781 86175
rect 219809 86147 219843 86175
rect 219871 86147 219919 86175
rect 219609 86113 219919 86147
rect 219609 86085 219657 86113
rect 219685 86085 219719 86113
rect 219747 86085 219781 86113
rect 219809 86085 219843 86113
rect 219871 86085 219919 86113
rect 219609 86051 219919 86085
rect 219609 86023 219657 86051
rect 219685 86023 219719 86051
rect 219747 86023 219781 86051
rect 219809 86023 219843 86051
rect 219871 86023 219919 86051
rect 219609 85989 219919 86023
rect 219609 85961 219657 85989
rect 219685 85961 219719 85989
rect 219747 85961 219781 85989
rect 219809 85961 219843 85989
rect 219871 85961 219919 85989
rect 219609 77175 219919 85961
rect 219609 77147 219657 77175
rect 219685 77147 219719 77175
rect 219747 77147 219781 77175
rect 219809 77147 219843 77175
rect 219871 77147 219919 77175
rect 219609 77113 219919 77147
rect 219609 77085 219657 77113
rect 219685 77085 219719 77113
rect 219747 77085 219781 77113
rect 219809 77085 219843 77113
rect 219871 77085 219919 77113
rect 219609 77051 219919 77085
rect 219609 77023 219657 77051
rect 219685 77023 219719 77051
rect 219747 77023 219781 77051
rect 219809 77023 219843 77051
rect 219871 77023 219919 77051
rect 219609 76989 219919 77023
rect 219609 76961 219657 76989
rect 219685 76961 219719 76989
rect 219747 76961 219781 76989
rect 219809 76961 219843 76989
rect 219871 76961 219919 76989
rect 219609 68175 219919 76961
rect 219609 68147 219657 68175
rect 219685 68147 219719 68175
rect 219747 68147 219781 68175
rect 219809 68147 219843 68175
rect 219871 68147 219919 68175
rect 219609 68113 219919 68147
rect 219609 68085 219657 68113
rect 219685 68085 219719 68113
rect 219747 68085 219781 68113
rect 219809 68085 219843 68113
rect 219871 68085 219919 68113
rect 219609 68051 219919 68085
rect 219609 68023 219657 68051
rect 219685 68023 219719 68051
rect 219747 68023 219781 68051
rect 219809 68023 219843 68051
rect 219871 68023 219919 68051
rect 219609 67989 219919 68023
rect 219609 67961 219657 67989
rect 219685 67961 219719 67989
rect 219747 67961 219781 67989
rect 219809 67961 219843 67989
rect 219871 67961 219919 67989
rect 219609 59175 219919 67961
rect 219609 59147 219657 59175
rect 219685 59147 219719 59175
rect 219747 59147 219781 59175
rect 219809 59147 219843 59175
rect 219871 59147 219919 59175
rect 219609 59113 219919 59147
rect 219609 59085 219657 59113
rect 219685 59085 219719 59113
rect 219747 59085 219781 59113
rect 219809 59085 219843 59113
rect 219871 59085 219919 59113
rect 219609 59051 219919 59085
rect 219609 59023 219657 59051
rect 219685 59023 219719 59051
rect 219747 59023 219781 59051
rect 219809 59023 219843 59051
rect 219871 59023 219919 59051
rect 219609 58989 219919 59023
rect 219609 58961 219657 58989
rect 219685 58961 219719 58989
rect 219747 58961 219781 58989
rect 219809 58961 219843 58989
rect 219871 58961 219919 58989
rect 219609 50175 219919 58961
rect 219609 50147 219657 50175
rect 219685 50147 219719 50175
rect 219747 50147 219781 50175
rect 219809 50147 219843 50175
rect 219871 50147 219919 50175
rect 219609 50113 219919 50147
rect 219609 50085 219657 50113
rect 219685 50085 219719 50113
rect 219747 50085 219781 50113
rect 219809 50085 219843 50113
rect 219871 50085 219919 50113
rect 219609 50051 219919 50085
rect 219609 50023 219657 50051
rect 219685 50023 219719 50051
rect 219747 50023 219781 50051
rect 219809 50023 219843 50051
rect 219871 50023 219919 50051
rect 219609 49989 219919 50023
rect 219609 49961 219657 49989
rect 219685 49961 219719 49989
rect 219747 49961 219781 49989
rect 219809 49961 219843 49989
rect 219871 49961 219919 49989
rect 219609 41175 219919 49961
rect 219609 41147 219657 41175
rect 219685 41147 219719 41175
rect 219747 41147 219781 41175
rect 219809 41147 219843 41175
rect 219871 41147 219919 41175
rect 219609 41113 219919 41147
rect 219609 41085 219657 41113
rect 219685 41085 219719 41113
rect 219747 41085 219781 41113
rect 219809 41085 219843 41113
rect 219871 41085 219919 41113
rect 219609 41051 219919 41085
rect 219609 41023 219657 41051
rect 219685 41023 219719 41051
rect 219747 41023 219781 41051
rect 219809 41023 219843 41051
rect 219871 41023 219919 41051
rect 219609 40989 219919 41023
rect 219609 40961 219657 40989
rect 219685 40961 219719 40989
rect 219747 40961 219781 40989
rect 219809 40961 219843 40989
rect 219871 40961 219919 40989
rect 219609 32175 219919 40961
rect 219609 32147 219657 32175
rect 219685 32147 219719 32175
rect 219747 32147 219781 32175
rect 219809 32147 219843 32175
rect 219871 32147 219919 32175
rect 219609 32113 219919 32147
rect 219609 32085 219657 32113
rect 219685 32085 219719 32113
rect 219747 32085 219781 32113
rect 219809 32085 219843 32113
rect 219871 32085 219919 32113
rect 219609 32051 219919 32085
rect 219609 32023 219657 32051
rect 219685 32023 219719 32051
rect 219747 32023 219781 32051
rect 219809 32023 219843 32051
rect 219871 32023 219919 32051
rect 219609 31989 219919 32023
rect 219609 31961 219657 31989
rect 219685 31961 219719 31989
rect 219747 31961 219781 31989
rect 219809 31961 219843 31989
rect 219871 31961 219919 31989
rect 219609 23175 219919 31961
rect 219609 23147 219657 23175
rect 219685 23147 219719 23175
rect 219747 23147 219781 23175
rect 219809 23147 219843 23175
rect 219871 23147 219919 23175
rect 219609 23113 219919 23147
rect 219609 23085 219657 23113
rect 219685 23085 219719 23113
rect 219747 23085 219781 23113
rect 219809 23085 219843 23113
rect 219871 23085 219919 23113
rect 219609 23051 219919 23085
rect 219609 23023 219657 23051
rect 219685 23023 219719 23051
rect 219747 23023 219781 23051
rect 219809 23023 219843 23051
rect 219871 23023 219919 23051
rect 219609 22989 219919 23023
rect 219609 22961 219657 22989
rect 219685 22961 219719 22989
rect 219747 22961 219781 22989
rect 219809 22961 219843 22989
rect 219871 22961 219919 22989
rect 219609 14175 219919 22961
rect 219609 14147 219657 14175
rect 219685 14147 219719 14175
rect 219747 14147 219781 14175
rect 219809 14147 219843 14175
rect 219871 14147 219919 14175
rect 219609 14113 219919 14147
rect 219609 14085 219657 14113
rect 219685 14085 219719 14113
rect 219747 14085 219781 14113
rect 219809 14085 219843 14113
rect 219871 14085 219919 14113
rect 219609 14051 219919 14085
rect 219609 14023 219657 14051
rect 219685 14023 219719 14051
rect 219747 14023 219781 14051
rect 219809 14023 219843 14051
rect 219871 14023 219919 14051
rect 219609 13989 219919 14023
rect 219609 13961 219657 13989
rect 219685 13961 219719 13989
rect 219747 13961 219781 13989
rect 219809 13961 219843 13989
rect 219871 13961 219919 13989
rect 219609 5175 219919 13961
rect 219609 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 219919 5175
rect 219609 5113 219919 5147
rect 219609 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 219919 5113
rect 219609 5051 219919 5085
rect 219609 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 219919 5051
rect 219609 4989 219919 5023
rect 219609 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 219919 4989
rect 219609 -560 219919 4961
rect 219609 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 219919 -560
rect 219609 -622 219919 -588
rect 219609 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 219919 -622
rect 219609 -684 219919 -650
rect 219609 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 219919 -684
rect 219609 -746 219919 -712
rect 219609 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 219919 -746
rect 219609 -822 219919 -774
rect 233109 92175 233419 100689
rect 233109 92147 233157 92175
rect 233185 92147 233219 92175
rect 233247 92147 233281 92175
rect 233309 92147 233343 92175
rect 233371 92147 233419 92175
rect 233109 92113 233419 92147
rect 233109 92085 233157 92113
rect 233185 92085 233219 92113
rect 233247 92085 233281 92113
rect 233309 92085 233343 92113
rect 233371 92085 233419 92113
rect 233109 92051 233419 92085
rect 233109 92023 233157 92051
rect 233185 92023 233219 92051
rect 233247 92023 233281 92051
rect 233309 92023 233343 92051
rect 233371 92023 233419 92051
rect 233109 91989 233419 92023
rect 233109 91961 233157 91989
rect 233185 91961 233219 91989
rect 233247 91961 233281 91989
rect 233309 91961 233343 91989
rect 233371 91961 233419 91989
rect 233109 83175 233419 91961
rect 233109 83147 233157 83175
rect 233185 83147 233219 83175
rect 233247 83147 233281 83175
rect 233309 83147 233343 83175
rect 233371 83147 233419 83175
rect 233109 83113 233419 83147
rect 233109 83085 233157 83113
rect 233185 83085 233219 83113
rect 233247 83085 233281 83113
rect 233309 83085 233343 83113
rect 233371 83085 233419 83113
rect 233109 83051 233419 83085
rect 233109 83023 233157 83051
rect 233185 83023 233219 83051
rect 233247 83023 233281 83051
rect 233309 83023 233343 83051
rect 233371 83023 233419 83051
rect 233109 82989 233419 83023
rect 233109 82961 233157 82989
rect 233185 82961 233219 82989
rect 233247 82961 233281 82989
rect 233309 82961 233343 82989
rect 233371 82961 233419 82989
rect 233109 74175 233419 82961
rect 233109 74147 233157 74175
rect 233185 74147 233219 74175
rect 233247 74147 233281 74175
rect 233309 74147 233343 74175
rect 233371 74147 233419 74175
rect 233109 74113 233419 74147
rect 233109 74085 233157 74113
rect 233185 74085 233219 74113
rect 233247 74085 233281 74113
rect 233309 74085 233343 74113
rect 233371 74085 233419 74113
rect 233109 74051 233419 74085
rect 233109 74023 233157 74051
rect 233185 74023 233219 74051
rect 233247 74023 233281 74051
rect 233309 74023 233343 74051
rect 233371 74023 233419 74051
rect 233109 73989 233419 74023
rect 233109 73961 233157 73989
rect 233185 73961 233219 73989
rect 233247 73961 233281 73989
rect 233309 73961 233343 73989
rect 233371 73961 233419 73989
rect 233109 65175 233419 73961
rect 233109 65147 233157 65175
rect 233185 65147 233219 65175
rect 233247 65147 233281 65175
rect 233309 65147 233343 65175
rect 233371 65147 233419 65175
rect 233109 65113 233419 65147
rect 233109 65085 233157 65113
rect 233185 65085 233219 65113
rect 233247 65085 233281 65113
rect 233309 65085 233343 65113
rect 233371 65085 233419 65113
rect 233109 65051 233419 65085
rect 233109 65023 233157 65051
rect 233185 65023 233219 65051
rect 233247 65023 233281 65051
rect 233309 65023 233343 65051
rect 233371 65023 233419 65051
rect 233109 64989 233419 65023
rect 233109 64961 233157 64989
rect 233185 64961 233219 64989
rect 233247 64961 233281 64989
rect 233309 64961 233343 64989
rect 233371 64961 233419 64989
rect 233109 56175 233419 64961
rect 233109 56147 233157 56175
rect 233185 56147 233219 56175
rect 233247 56147 233281 56175
rect 233309 56147 233343 56175
rect 233371 56147 233419 56175
rect 233109 56113 233419 56147
rect 233109 56085 233157 56113
rect 233185 56085 233219 56113
rect 233247 56085 233281 56113
rect 233309 56085 233343 56113
rect 233371 56085 233419 56113
rect 233109 56051 233419 56085
rect 233109 56023 233157 56051
rect 233185 56023 233219 56051
rect 233247 56023 233281 56051
rect 233309 56023 233343 56051
rect 233371 56023 233419 56051
rect 233109 55989 233419 56023
rect 233109 55961 233157 55989
rect 233185 55961 233219 55989
rect 233247 55961 233281 55989
rect 233309 55961 233343 55989
rect 233371 55961 233419 55989
rect 233109 47175 233419 55961
rect 233109 47147 233157 47175
rect 233185 47147 233219 47175
rect 233247 47147 233281 47175
rect 233309 47147 233343 47175
rect 233371 47147 233419 47175
rect 233109 47113 233419 47147
rect 233109 47085 233157 47113
rect 233185 47085 233219 47113
rect 233247 47085 233281 47113
rect 233309 47085 233343 47113
rect 233371 47085 233419 47113
rect 233109 47051 233419 47085
rect 233109 47023 233157 47051
rect 233185 47023 233219 47051
rect 233247 47023 233281 47051
rect 233309 47023 233343 47051
rect 233371 47023 233419 47051
rect 233109 46989 233419 47023
rect 233109 46961 233157 46989
rect 233185 46961 233219 46989
rect 233247 46961 233281 46989
rect 233309 46961 233343 46989
rect 233371 46961 233419 46989
rect 233109 38175 233419 46961
rect 233109 38147 233157 38175
rect 233185 38147 233219 38175
rect 233247 38147 233281 38175
rect 233309 38147 233343 38175
rect 233371 38147 233419 38175
rect 233109 38113 233419 38147
rect 233109 38085 233157 38113
rect 233185 38085 233219 38113
rect 233247 38085 233281 38113
rect 233309 38085 233343 38113
rect 233371 38085 233419 38113
rect 233109 38051 233419 38085
rect 233109 38023 233157 38051
rect 233185 38023 233219 38051
rect 233247 38023 233281 38051
rect 233309 38023 233343 38051
rect 233371 38023 233419 38051
rect 233109 37989 233419 38023
rect 233109 37961 233157 37989
rect 233185 37961 233219 37989
rect 233247 37961 233281 37989
rect 233309 37961 233343 37989
rect 233371 37961 233419 37989
rect 233109 29175 233419 37961
rect 233109 29147 233157 29175
rect 233185 29147 233219 29175
rect 233247 29147 233281 29175
rect 233309 29147 233343 29175
rect 233371 29147 233419 29175
rect 233109 29113 233419 29147
rect 233109 29085 233157 29113
rect 233185 29085 233219 29113
rect 233247 29085 233281 29113
rect 233309 29085 233343 29113
rect 233371 29085 233419 29113
rect 233109 29051 233419 29085
rect 233109 29023 233157 29051
rect 233185 29023 233219 29051
rect 233247 29023 233281 29051
rect 233309 29023 233343 29051
rect 233371 29023 233419 29051
rect 233109 28989 233419 29023
rect 233109 28961 233157 28989
rect 233185 28961 233219 28989
rect 233247 28961 233281 28989
rect 233309 28961 233343 28989
rect 233371 28961 233419 28989
rect 233109 20175 233419 28961
rect 233109 20147 233157 20175
rect 233185 20147 233219 20175
rect 233247 20147 233281 20175
rect 233309 20147 233343 20175
rect 233371 20147 233419 20175
rect 233109 20113 233419 20147
rect 233109 20085 233157 20113
rect 233185 20085 233219 20113
rect 233247 20085 233281 20113
rect 233309 20085 233343 20113
rect 233371 20085 233419 20113
rect 233109 20051 233419 20085
rect 233109 20023 233157 20051
rect 233185 20023 233219 20051
rect 233247 20023 233281 20051
rect 233309 20023 233343 20051
rect 233371 20023 233419 20051
rect 233109 19989 233419 20023
rect 233109 19961 233157 19989
rect 233185 19961 233219 19989
rect 233247 19961 233281 19989
rect 233309 19961 233343 19989
rect 233371 19961 233419 19989
rect 233109 11175 233419 19961
rect 233109 11147 233157 11175
rect 233185 11147 233219 11175
rect 233247 11147 233281 11175
rect 233309 11147 233343 11175
rect 233371 11147 233419 11175
rect 233109 11113 233419 11147
rect 233109 11085 233157 11113
rect 233185 11085 233219 11113
rect 233247 11085 233281 11113
rect 233309 11085 233343 11113
rect 233371 11085 233419 11113
rect 233109 11051 233419 11085
rect 233109 11023 233157 11051
rect 233185 11023 233219 11051
rect 233247 11023 233281 11051
rect 233309 11023 233343 11051
rect 233371 11023 233419 11051
rect 233109 10989 233419 11023
rect 233109 10961 233157 10989
rect 233185 10961 233219 10989
rect 233247 10961 233281 10989
rect 233309 10961 233343 10989
rect 233371 10961 233419 10989
rect 233109 2175 233419 10961
rect 233109 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 233419 2175
rect 233109 2113 233419 2147
rect 233109 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 233419 2113
rect 233109 2051 233419 2085
rect 233109 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 233419 2051
rect 233109 1989 233419 2023
rect 233109 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 233419 1989
rect 233109 -80 233419 1961
rect 233109 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 233419 -80
rect 233109 -142 233419 -108
rect 233109 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 233419 -142
rect 233109 -204 233419 -170
rect 233109 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 233419 -204
rect 233109 -266 233419 -232
rect 233109 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 233419 -266
rect 233109 -822 233419 -294
rect 234969 95175 235279 100689
rect 234969 95147 235017 95175
rect 235045 95147 235079 95175
rect 235107 95147 235141 95175
rect 235169 95147 235203 95175
rect 235231 95147 235279 95175
rect 234969 95113 235279 95147
rect 234969 95085 235017 95113
rect 235045 95085 235079 95113
rect 235107 95085 235141 95113
rect 235169 95085 235203 95113
rect 235231 95085 235279 95113
rect 234969 95051 235279 95085
rect 234969 95023 235017 95051
rect 235045 95023 235079 95051
rect 235107 95023 235141 95051
rect 235169 95023 235203 95051
rect 235231 95023 235279 95051
rect 234969 94989 235279 95023
rect 234969 94961 235017 94989
rect 235045 94961 235079 94989
rect 235107 94961 235141 94989
rect 235169 94961 235203 94989
rect 235231 94961 235279 94989
rect 234969 86175 235279 94961
rect 234969 86147 235017 86175
rect 235045 86147 235079 86175
rect 235107 86147 235141 86175
rect 235169 86147 235203 86175
rect 235231 86147 235279 86175
rect 234969 86113 235279 86147
rect 234969 86085 235017 86113
rect 235045 86085 235079 86113
rect 235107 86085 235141 86113
rect 235169 86085 235203 86113
rect 235231 86085 235279 86113
rect 234969 86051 235279 86085
rect 234969 86023 235017 86051
rect 235045 86023 235079 86051
rect 235107 86023 235141 86051
rect 235169 86023 235203 86051
rect 235231 86023 235279 86051
rect 234969 85989 235279 86023
rect 234969 85961 235017 85989
rect 235045 85961 235079 85989
rect 235107 85961 235141 85989
rect 235169 85961 235203 85989
rect 235231 85961 235279 85989
rect 234969 77175 235279 85961
rect 234969 77147 235017 77175
rect 235045 77147 235079 77175
rect 235107 77147 235141 77175
rect 235169 77147 235203 77175
rect 235231 77147 235279 77175
rect 234969 77113 235279 77147
rect 234969 77085 235017 77113
rect 235045 77085 235079 77113
rect 235107 77085 235141 77113
rect 235169 77085 235203 77113
rect 235231 77085 235279 77113
rect 234969 77051 235279 77085
rect 234969 77023 235017 77051
rect 235045 77023 235079 77051
rect 235107 77023 235141 77051
rect 235169 77023 235203 77051
rect 235231 77023 235279 77051
rect 234969 76989 235279 77023
rect 234969 76961 235017 76989
rect 235045 76961 235079 76989
rect 235107 76961 235141 76989
rect 235169 76961 235203 76989
rect 235231 76961 235279 76989
rect 234969 68175 235279 76961
rect 234969 68147 235017 68175
rect 235045 68147 235079 68175
rect 235107 68147 235141 68175
rect 235169 68147 235203 68175
rect 235231 68147 235279 68175
rect 234969 68113 235279 68147
rect 234969 68085 235017 68113
rect 235045 68085 235079 68113
rect 235107 68085 235141 68113
rect 235169 68085 235203 68113
rect 235231 68085 235279 68113
rect 234969 68051 235279 68085
rect 234969 68023 235017 68051
rect 235045 68023 235079 68051
rect 235107 68023 235141 68051
rect 235169 68023 235203 68051
rect 235231 68023 235279 68051
rect 234969 67989 235279 68023
rect 234969 67961 235017 67989
rect 235045 67961 235079 67989
rect 235107 67961 235141 67989
rect 235169 67961 235203 67989
rect 235231 67961 235279 67989
rect 234969 59175 235279 67961
rect 234969 59147 235017 59175
rect 235045 59147 235079 59175
rect 235107 59147 235141 59175
rect 235169 59147 235203 59175
rect 235231 59147 235279 59175
rect 234969 59113 235279 59147
rect 234969 59085 235017 59113
rect 235045 59085 235079 59113
rect 235107 59085 235141 59113
rect 235169 59085 235203 59113
rect 235231 59085 235279 59113
rect 234969 59051 235279 59085
rect 234969 59023 235017 59051
rect 235045 59023 235079 59051
rect 235107 59023 235141 59051
rect 235169 59023 235203 59051
rect 235231 59023 235279 59051
rect 234969 58989 235279 59023
rect 234969 58961 235017 58989
rect 235045 58961 235079 58989
rect 235107 58961 235141 58989
rect 235169 58961 235203 58989
rect 235231 58961 235279 58989
rect 234969 50175 235279 58961
rect 234969 50147 235017 50175
rect 235045 50147 235079 50175
rect 235107 50147 235141 50175
rect 235169 50147 235203 50175
rect 235231 50147 235279 50175
rect 234969 50113 235279 50147
rect 234969 50085 235017 50113
rect 235045 50085 235079 50113
rect 235107 50085 235141 50113
rect 235169 50085 235203 50113
rect 235231 50085 235279 50113
rect 234969 50051 235279 50085
rect 234969 50023 235017 50051
rect 235045 50023 235079 50051
rect 235107 50023 235141 50051
rect 235169 50023 235203 50051
rect 235231 50023 235279 50051
rect 234969 49989 235279 50023
rect 234969 49961 235017 49989
rect 235045 49961 235079 49989
rect 235107 49961 235141 49989
rect 235169 49961 235203 49989
rect 235231 49961 235279 49989
rect 234969 41175 235279 49961
rect 234969 41147 235017 41175
rect 235045 41147 235079 41175
rect 235107 41147 235141 41175
rect 235169 41147 235203 41175
rect 235231 41147 235279 41175
rect 234969 41113 235279 41147
rect 234969 41085 235017 41113
rect 235045 41085 235079 41113
rect 235107 41085 235141 41113
rect 235169 41085 235203 41113
rect 235231 41085 235279 41113
rect 234969 41051 235279 41085
rect 234969 41023 235017 41051
rect 235045 41023 235079 41051
rect 235107 41023 235141 41051
rect 235169 41023 235203 41051
rect 235231 41023 235279 41051
rect 234969 40989 235279 41023
rect 234969 40961 235017 40989
rect 235045 40961 235079 40989
rect 235107 40961 235141 40989
rect 235169 40961 235203 40989
rect 235231 40961 235279 40989
rect 234969 32175 235279 40961
rect 234969 32147 235017 32175
rect 235045 32147 235079 32175
rect 235107 32147 235141 32175
rect 235169 32147 235203 32175
rect 235231 32147 235279 32175
rect 234969 32113 235279 32147
rect 234969 32085 235017 32113
rect 235045 32085 235079 32113
rect 235107 32085 235141 32113
rect 235169 32085 235203 32113
rect 235231 32085 235279 32113
rect 234969 32051 235279 32085
rect 234969 32023 235017 32051
rect 235045 32023 235079 32051
rect 235107 32023 235141 32051
rect 235169 32023 235203 32051
rect 235231 32023 235279 32051
rect 234969 31989 235279 32023
rect 234969 31961 235017 31989
rect 235045 31961 235079 31989
rect 235107 31961 235141 31989
rect 235169 31961 235203 31989
rect 235231 31961 235279 31989
rect 234969 23175 235279 31961
rect 234969 23147 235017 23175
rect 235045 23147 235079 23175
rect 235107 23147 235141 23175
rect 235169 23147 235203 23175
rect 235231 23147 235279 23175
rect 234969 23113 235279 23147
rect 234969 23085 235017 23113
rect 235045 23085 235079 23113
rect 235107 23085 235141 23113
rect 235169 23085 235203 23113
rect 235231 23085 235279 23113
rect 234969 23051 235279 23085
rect 234969 23023 235017 23051
rect 235045 23023 235079 23051
rect 235107 23023 235141 23051
rect 235169 23023 235203 23051
rect 235231 23023 235279 23051
rect 234969 22989 235279 23023
rect 234969 22961 235017 22989
rect 235045 22961 235079 22989
rect 235107 22961 235141 22989
rect 235169 22961 235203 22989
rect 235231 22961 235279 22989
rect 234969 14175 235279 22961
rect 234969 14147 235017 14175
rect 235045 14147 235079 14175
rect 235107 14147 235141 14175
rect 235169 14147 235203 14175
rect 235231 14147 235279 14175
rect 234969 14113 235279 14147
rect 234969 14085 235017 14113
rect 235045 14085 235079 14113
rect 235107 14085 235141 14113
rect 235169 14085 235203 14113
rect 235231 14085 235279 14113
rect 234969 14051 235279 14085
rect 234969 14023 235017 14051
rect 235045 14023 235079 14051
rect 235107 14023 235141 14051
rect 235169 14023 235203 14051
rect 235231 14023 235279 14051
rect 234969 13989 235279 14023
rect 234969 13961 235017 13989
rect 235045 13961 235079 13989
rect 235107 13961 235141 13989
rect 235169 13961 235203 13989
rect 235231 13961 235279 13989
rect 234969 5175 235279 13961
rect 234969 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 235279 5175
rect 234969 5113 235279 5147
rect 234969 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 235279 5113
rect 234969 5051 235279 5085
rect 234969 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 235279 5051
rect 234969 4989 235279 5023
rect 234969 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 235279 4989
rect 234969 -560 235279 4961
rect 234969 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 235279 -560
rect 234969 -622 235279 -588
rect 234969 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 235279 -622
rect 234969 -684 235279 -650
rect 234969 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 235279 -684
rect 234969 -746 235279 -712
rect 234969 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 235279 -746
rect 234969 -822 235279 -774
rect 248469 92175 248779 100689
rect 248469 92147 248517 92175
rect 248545 92147 248579 92175
rect 248607 92147 248641 92175
rect 248669 92147 248703 92175
rect 248731 92147 248779 92175
rect 248469 92113 248779 92147
rect 248469 92085 248517 92113
rect 248545 92085 248579 92113
rect 248607 92085 248641 92113
rect 248669 92085 248703 92113
rect 248731 92085 248779 92113
rect 248469 92051 248779 92085
rect 248469 92023 248517 92051
rect 248545 92023 248579 92051
rect 248607 92023 248641 92051
rect 248669 92023 248703 92051
rect 248731 92023 248779 92051
rect 248469 91989 248779 92023
rect 248469 91961 248517 91989
rect 248545 91961 248579 91989
rect 248607 91961 248641 91989
rect 248669 91961 248703 91989
rect 248731 91961 248779 91989
rect 248469 83175 248779 91961
rect 248469 83147 248517 83175
rect 248545 83147 248579 83175
rect 248607 83147 248641 83175
rect 248669 83147 248703 83175
rect 248731 83147 248779 83175
rect 248469 83113 248779 83147
rect 248469 83085 248517 83113
rect 248545 83085 248579 83113
rect 248607 83085 248641 83113
rect 248669 83085 248703 83113
rect 248731 83085 248779 83113
rect 248469 83051 248779 83085
rect 248469 83023 248517 83051
rect 248545 83023 248579 83051
rect 248607 83023 248641 83051
rect 248669 83023 248703 83051
rect 248731 83023 248779 83051
rect 248469 82989 248779 83023
rect 248469 82961 248517 82989
rect 248545 82961 248579 82989
rect 248607 82961 248641 82989
rect 248669 82961 248703 82989
rect 248731 82961 248779 82989
rect 248469 74175 248779 82961
rect 248469 74147 248517 74175
rect 248545 74147 248579 74175
rect 248607 74147 248641 74175
rect 248669 74147 248703 74175
rect 248731 74147 248779 74175
rect 248469 74113 248779 74147
rect 248469 74085 248517 74113
rect 248545 74085 248579 74113
rect 248607 74085 248641 74113
rect 248669 74085 248703 74113
rect 248731 74085 248779 74113
rect 248469 74051 248779 74085
rect 248469 74023 248517 74051
rect 248545 74023 248579 74051
rect 248607 74023 248641 74051
rect 248669 74023 248703 74051
rect 248731 74023 248779 74051
rect 248469 73989 248779 74023
rect 248469 73961 248517 73989
rect 248545 73961 248579 73989
rect 248607 73961 248641 73989
rect 248669 73961 248703 73989
rect 248731 73961 248779 73989
rect 248469 65175 248779 73961
rect 248469 65147 248517 65175
rect 248545 65147 248579 65175
rect 248607 65147 248641 65175
rect 248669 65147 248703 65175
rect 248731 65147 248779 65175
rect 248469 65113 248779 65147
rect 248469 65085 248517 65113
rect 248545 65085 248579 65113
rect 248607 65085 248641 65113
rect 248669 65085 248703 65113
rect 248731 65085 248779 65113
rect 248469 65051 248779 65085
rect 248469 65023 248517 65051
rect 248545 65023 248579 65051
rect 248607 65023 248641 65051
rect 248669 65023 248703 65051
rect 248731 65023 248779 65051
rect 248469 64989 248779 65023
rect 248469 64961 248517 64989
rect 248545 64961 248579 64989
rect 248607 64961 248641 64989
rect 248669 64961 248703 64989
rect 248731 64961 248779 64989
rect 248469 56175 248779 64961
rect 248469 56147 248517 56175
rect 248545 56147 248579 56175
rect 248607 56147 248641 56175
rect 248669 56147 248703 56175
rect 248731 56147 248779 56175
rect 248469 56113 248779 56147
rect 248469 56085 248517 56113
rect 248545 56085 248579 56113
rect 248607 56085 248641 56113
rect 248669 56085 248703 56113
rect 248731 56085 248779 56113
rect 248469 56051 248779 56085
rect 248469 56023 248517 56051
rect 248545 56023 248579 56051
rect 248607 56023 248641 56051
rect 248669 56023 248703 56051
rect 248731 56023 248779 56051
rect 248469 55989 248779 56023
rect 248469 55961 248517 55989
rect 248545 55961 248579 55989
rect 248607 55961 248641 55989
rect 248669 55961 248703 55989
rect 248731 55961 248779 55989
rect 248469 47175 248779 55961
rect 248469 47147 248517 47175
rect 248545 47147 248579 47175
rect 248607 47147 248641 47175
rect 248669 47147 248703 47175
rect 248731 47147 248779 47175
rect 248469 47113 248779 47147
rect 248469 47085 248517 47113
rect 248545 47085 248579 47113
rect 248607 47085 248641 47113
rect 248669 47085 248703 47113
rect 248731 47085 248779 47113
rect 248469 47051 248779 47085
rect 248469 47023 248517 47051
rect 248545 47023 248579 47051
rect 248607 47023 248641 47051
rect 248669 47023 248703 47051
rect 248731 47023 248779 47051
rect 248469 46989 248779 47023
rect 248469 46961 248517 46989
rect 248545 46961 248579 46989
rect 248607 46961 248641 46989
rect 248669 46961 248703 46989
rect 248731 46961 248779 46989
rect 248469 38175 248779 46961
rect 248469 38147 248517 38175
rect 248545 38147 248579 38175
rect 248607 38147 248641 38175
rect 248669 38147 248703 38175
rect 248731 38147 248779 38175
rect 248469 38113 248779 38147
rect 248469 38085 248517 38113
rect 248545 38085 248579 38113
rect 248607 38085 248641 38113
rect 248669 38085 248703 38113
rect 248731 38085 248779 38113
rect 248469 38051 248779 38085
rect 248469 38023 248517 38051
rect 248545 38023 248579 38051
rect 248607 38023 248641 38051
rect 248669 38023 248703 38051
rect 248731 38023 248779 38051
rect 248469 37989 248779 38023
rect 248469 37961 248517 37989
rect 248545 37961 248579 37989
rect 248607 37961 248641 37989
rect 248669 37961 248703 37989
rect 248731 37961 248779 37989
rect 248469 29175 248779 37961
rect 248469 29147 248517 29175
rect 248545 29147 248579 29175
rect 248607 29147 248641 29175
rect 248669 29147 248703 29175
rect 248731 29147 248779 29175
rect 248469 29113 248779 29147
rect 248469 29085 248517 29113
rect 248545 29085 248579 29113
rect 248607 29085 248641 29113
rect 248669 29085 248703 29113
rect 248731 29085 248779 29113
rect 248469 29051 248779 29085
rect 248469 29023 248517 29051
rect 248545 29023 248579 29051
rect 248607 29023 248641 29051
rect 248669 29023 248703 29051
rect 248731 29023 248779 29051
rect 248469 28989 248779 29023
rect 248469 28961 248517 28989
rect 248545 28961 248579 28989
rect 248607 28961 248641 28989
rect 248669 28961 248703 28989
rect 248731 28961 248779 28989
rect 248469 20175 248779 28961
rect 248469 20147 248517 20175
rect 248545 20147 248579 20175
rect 248607 20147 248641 20175
rect 248669 20147 248703 20175
rect 248731 20147 248779 20175
rect 248469 20113 248779 20147
rect 248469 20085 248517 20113
rect 248545 20085 248579 20113
rect 248607 20085 248641 20113
rect 248669 20085 248703 20113
rect 248731 20085 248779 20113
rect 248469 20051 248779 20085
rect 248469 20023 248517 20051
rect 248545 20023 248579 20051
rect 248607 20023 248641 20051
rect 248669 20023 248703 20051
rect 248731 20023 248779 20051
rect 248469 19989 248779 20023
rect 248469 19961 248517 19989
rect 248545 19961 248579 19989
rect 248607 19961 248641 19989
rect 248669 19961 248703 19989
rect 248731 19961 248779 19989
rect 248469 11175 248779 19961
rect 248469 11147 248517 11175
rect 248545 11147 248579 11175
rect 248607 11147 248641 11175
rect 248669 11147 248703 11175
rect 248731 11147 248779 11175
rect 248469 11113 248779 11147
rect 248469 11085 248517 11113
rect 248545 11085 248579 11113
rect 248607 11085 248641 11113
rect 248669 11085 248703 11113
rect 248731 11085 248779 11113
rect 248469 11051 248779 11085
rect 248469 11023 248517 11051
rect 248545 11023 248579 11051
rect 248607 11023 248641 11051
rect 248669 11023 248703 11051
rect 248731 11023 248779 11051
rect 248469 10989 248779 11023
rect 248469 10961 248517 10989
rect 248545 10961 248579 10989
rect 248607 10961 248641 10989
rect 248669 10961 248703 10989
rect 248731 10961 248779 10989
rect 248469 2175 248779 10961
rect 248469 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 248779 2175
rect 248469 2113 248779 2147
rect 248469 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 248779 2113
rect 248469 2051 248779 2085
rect 248469 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 248779 2051
rect 248469 1989 248779 2023
rect 248469 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 248779 1989
rect 248469 -80 248779 1961
rect 248469 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 248779 -80
rect 248469 -142 248779 -108
rect 248469 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 248779 -142
rect 248469 -204 248779 -170
rect 248469 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 248779 -204
rect 248469 -266 248779 -232
rect 248469 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 248779 -266
rect 248469 -822 248779 -294
rect 250329 95175 250639 100689
rect 250329 95147 250377 95175
rect 250405 95147 250439 95175
rect 250467 95147 250501 95175
rect 250529 95147 250563 95175
rect 250591 95147 250639 95175
rect 250329 95113 250639 95147
rect 250329 95085 250377 95113
rect 250405 95085 250439 95113
rect 250467 95085 250501 95113
rect 250529 95085 250563 95113
rect 250591 95085 250639 95113
rect 250329 95051 250639 95085
rect 250329 95023 250377 95051
rect 250405 95023 250439 95051
rect 250467 95023 250501 95051
rect 250529 95023 250563 95051
rect 250591 95023 250639 95051
rect 250329 94989 250639 95023
rect 250329 94961 250377 94989
rect 250405 94961 250439 94989
rect 250467 94961 250501 94989
rect 250529 94961 250563 94989
rect 250591 94961 250639 94989
rect 250329 86175 250639 94961
rect 250329 86147 250377 86175
rect 250405 86147 250439 86175
rect 250467 86147 250501 86175
rect 250529 86147 250563 86175
rect 250591 86147 250639 86175
rect 250329 86113 250639 86147
rect 250329 86085 250377 86113
rect 250405 86085 250439 86113
rect 250467 86085 250501 86113
rect 250529 86085 250563 86113
rect 250591 86085 250639 86113
rect 250329 86051 250639 86085
rect 250329 86023 250377 86051
rect 250405 86023 250439 86051
rect 250467 86023 250501 86051
rect 250529 86023 250563 86051
rect 250591 86023 250639 86051
rect 250329 85989 250639 86023
rect 250329 85961 250377 85989
rect 250405 85961 250439 85989
rect 250467 85961 250501 85989
rect 250529 85961 250563 85989
rect 250591 85961 250639 85989
rect 250329 77175 250639 85961
rect 250329 77147 250377 77175
rect 250405 77147 250439 77175
rect 250467 77147 250501 77175
rect 250529 77147 250563 77175
rect 250591 77147 250639 77175
rect 250329 77113 250639 77147
rect 250329 77085 250377 77113
rect 250405 77085 250439 77113
rect 250467 77085 250501 77113
rect 250529 77085 250563 77113
rect 250591 77085 250639 77113
rect 250329 77051 250639 77085
rect 250329 77023 250377 77051
rect 250405 77023 250439 77051
rect 250467 77023 250501 77051
rect 250529 77023 250563 77051
rect 250591 77023 250639 77051
rect 250329 76989 250639 77023
rect 250329 76961 250377 76989
rect 250405 76961 250439 76989
rect 250467 76961 250501 76989
rect 250529 76961 250563 76989
rect 250591 76961 250639 76989
rect 250329 68175 250639 76961
rect 250329 68147 250377 68175
rect 250405 68147 250439 68175
rect 250467 68147 250501 68175
rect 250529 68147 250563 68175
rect 250591 68147 250639 68175
rect 250329 68113 250639 68147
rect 250329 68085 250377 68113
rect 250405 68085 250439 68113
rect 250467 68085 250501 68113
rect 250529 68085 250563 68113
rect 250591 68085 250639 68113
rect 250329 68051 250639 68085
rect 250329 68023 250377 68051
rect 250405 68023 250439 68051
rect 250467 68023 250501 68051
rect 250529 68023 250563 68051
rect 250591 68023 250639 68051
rect 250329 67989 250639 68023
rect 250329 67961 250377 67989
rect 250405 67961 250439 67989
rect 250467 67961 250501 67989
rect 250529 67961 250563 67989
rect 250591 67961 250639 67989
rect 250329 59175 250639 67961
rect 250329 59147 250377 59175
rect 250405 59147 250439 59175
rect 250467 59147 250501 59175
rect 250529 59147 250563 59175
rect 250591 59147 250639 59175
rect 250329 59113 250639 59147
rect 250329 59085 250377 59113
rect 250405 59085 250439 59113
rect 250467 59085 250501 59113
rect 250529 59085 250563 59113
rect 250591 59085 250639 59113
rect 250329 59051 250639 59085
rect 250329 59023 250377 59051
rect 250405 59023 250439 59051
rect 250467 59023 250501 59051
rect 250529 59023 250563 59051
rect 250591 59023 250639 59051
rect 250329 58989 250639 59023
rect 250329 58961 250377 58989
rect 250405 58961 250439 58989
rect 250467 58961 250501 58989
rect 250529 58961 250563 58989
rect 250591 58961 250639 58989
rect 250329 50175 250639 58961
rect 250329 50147 250377 50175
rect 250405 50147 250439 50175
rect 250467 50147 250501 50175
rect 250529 50147 250563 50175
rect 250591 50147 250639 50175
rect 250329 50113 250639 50147
rect 250329 50085 250377 50113
rect 250405 50085 250439 50113
rect 250467 50085 250501 50113
rect 250529 50085 250563 50113
rect 250591 50085 250639 50113
rect 250329 50051 250639 50085
rect 250329 50023 250377 50051
rect 250405 50023 250439 50051
rect 250467 50023 250501 50051
rect 250529 50023 250563 50051
rect 250591 50023 250639 50051
rect 250329 49989 250639 50023
rect 250329 49961 250377 49989
rect 250405 49961 250439 49989
rect 250467 49961 250501 49989
rect 250529 49961 250563 49989
rect 250591 49961 250639 49989
rect 250329 41175 250639 49961
rect 250329 41147 250377 41175
rect 250405 41147 250439 41175
rect 250467 41147 250501 41175
rect 250529 41147 250563 41175
rect 250591 41147 250639 41175
rect 250329 41113 250639 41147
rect 250329 41085 250377 41113
rect 250405 41085 250439 41113
rect 250467 41085 250501 41113
rect 250529 41085 250563 41113
rect 250591 41085 250639 41113
rect 250329 41051 250639 41085
rect 250329 41023 250377 41051
rect 250405 41023 250439 41051
rect 250467 41023 250501 41051
rect 250529 41023 250563 41051
rect 250591 41023 250639 41051
rect 250329 40989 250639 41023
rect 250329 40961 250377 40989
rect 250405 40961 250439 40989
rect 250467 40961 250501 40989
rect 250529 40961 250563 40989
rect 250591 40961 250639 40989
rect 250329 32175 250639 40961
rect 250329 32147 250377 32175
rect 250405 32147 250439 32175
rect 250467 32147 250501 32175
rect 250529 32147 250563 32175
rect 250591 32147 250639 32175
rect 250329 32113 250639 32147
rect 250329 32085 250377 32113
rect 250405 32085 250439 32113
rect 250467 32085 250501 32113
rect 250529 32085 250563 32113
rect 250591 32085 250639 32113
rect 250329 32051 250639 32085
rect 250329 32023 250377 32051
rect 250405 32023 250439 32051
rect 250467 32023 250501 32051
rect 250529 32023 250563 32051
rect 250591 32023 250639 32051
rect 250329 31989 250639 32023
rect 250329 31961 250377 31989
rect 250405 31961 250439 31989
rect 250467 31961 250501 31989
rect 250529 31961 250563 31989
rect 250591 31961 250639 31989
rect 250329 23175 250639 31961
rect 250329 23147 250377 23175
rect 250405 23147 250439 23175
rect 250467 23147 250501 23175
rect 250529 23147 250563 23175
rect 250591 23147 250639 23175
rect 250329 23113 250639 23147
rect 250329 23085 250377 23113
rect 250405 23085 250439 23113
rect 250467 23085 250501 23113
rect 250529 23085 250563 23113
rect 250591 23085 250639 23113
rect 250329 23051 250639 23085
rect 250329 23023 250377 23051
rect 250405 23023 250439 23051
rect 250467 23023 250501 23051
rect 250529 23023 250563 23051
rect 250591 23023 250639 23051
rect 250329 22989 250639 23023
rect 250329 22961 250377 22989
rect 250405 22961 250439 22989
rect 250467 22961 250501 22989
rect 250529 22961 250563 22989
rect 250591 22961 250639 22989
rect 250329 14175 250639 22961
rect 250329 14147 250377 14175
rect 250405 14147 250439 14175
rect 250467 14147 250501 14175
rect 250529 14147 250563 14175
rect 250591 14147 250639 14175
rect 250329 14113 250639 14147
rect 250329 14085 250377 14113
rect 250405 14085 250439 14113
rect 250467 14085 250501 14113
rect 250529 14085 250563 14113
rect 250591 14085 250639 14113
rect 250329 14051 250639 14085
rect 250329 14023 250377 14051
rect 250405 14023 250439 14051
rect 250467 14023 250501 14051
rect 250529 14023 250563 14051
rect 250591 14023 250639 14051
rect 250329 13989 250639 14023
rect 250329 13961 250377 13989
rect 250405 13961 250439 13989
rect 250467 13961 250501 13989
rect 250529 13961 250563 13989
rect 250591 13961 250639 13989
rect 250329 5175 250639 13961
rect 250329 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 250639 5175
rect 250329 5113 250639 5147
rect 250329 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 250639 5113
rect 250329 5051 250639 5085
rect 250329 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 250639 5051
rect 250329 4989 250639 5023
rect 250329 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 250639 4989
rect 250329 -560 250639 4961
rect 250329 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 250639 -560
rect 250329 -622 250639 -588
rect 250329 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 250639 -622
rect 250329 -684 250639 -650
rect 250329 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 250639 -684
rect 250329 -746 250639 -712
rect 250329 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 250639 -746
rect 250329 -822 250639 -774
rect 263829 92175 264139 100689
rect 263829 92147 263877 92175
rect 263905 92147 263939 92175
rect 263967 92147 264001 92175
rect 264029 92147 264063 92175
rect 264091 92147 264139 92175
rect 263829 92113 264139 92147
rect 263829 92085 263877 92113
rect 263905 92085 263939 92113
rect 263967 92085 264001 92113
rect 264029 92085 264063 92113
rect 264091 92085 264139 92113
rect 263829 92051 264139 92085
rect 263829 92023 263877 92051
rect 263905 92023 263939 92051
rect 263967 92023 264001 92051
rect 264029 92023 264063 92051
rect 264091 92023 264139 92051
rect 263829 91989 264139 92023
rect 263829 91961 263877 91989
rect 263905 91961 263939 91989
rect 263967 91961 264001 91989
rect 264029 91961 264063 91989
rect 264091 91961 264139 91989
rect 263829 83175 264139 91961
rect 263829 83147 263877 83175
rect 263905 83147 263939 83175
rect 263967 83147 264001 83175
rect 264029 83147 264063 83175
rect 264091 83147 264139 83175
rect 263829 83113 264139 83147
rect 263829 83085 263877 83113
rect 263905 83085 263939 83113
rect 263967 83085 264001 83113
rect 264029 83085 264063 83113
rect 264091 83085 264139 83113
rect 263829 83051 264139 83085
rect 263829 83023 263877 83051
rect 263905 83023 263939 83051
rect 263967 83023 264001 83051
rect 264029 83023 264063 83051
rect 264091 83023 264139 83051
rect 263829 82989 264139 83023
rect 263829 82961 263877 82989
rect 263905 82961 263939 82989
rect 263967 82961 264001 82989
rect 264029 82961 264063 82989
rect 264091 82961 264139 82989
rect 263829 74175 264139 82961
rect 263829 74147 263877 74175
rect 263905 74147 263939 74175
rect 263967 74147 264001 74175
rect 264029 74147 264063 74175
rect 264091 74147 264139 74175
rect 263829 74113 264139 74147
rect 263829 74085 263877 74113
rect 263905 74085 263939 74113
rect 263967 74085 264001 74113
rect 264029 74085 264063 74113
rect 264091 74085 264139 74113
rect 263829 74051 264139 74085
rect 263829 74023 263877 74051
rect 263905 74023 263939 74051
rect 263967 74023 264001 74051
rect 264029 74023 264063 74051
rect 264091 74023 264139 74051
rect 263829 73989 264139 74023
rect 263829 73961 263877 73989
rect 263905 73961 263939 73989
rect 263967 73961 264001 73989
rect 264029 73961 264063 73989
rect 264091 73961 264139 73989
rect 263829 65175 264139 73961
rect 263829 65147 263877 65175
rect 263905 65147 263939 65175
rect 263967 65147 264001 65175
rect 264029 65147 264063 65175
rect 264091 65147 264139 65175
rect 263829 65113 264139 65147
rect 263829 65085 263877 65113
rect 263905 65085 263939 65113
rect 263967 65085 264001 65113
rect 264029 65085 264063 65113
rect 264091 65085 264139 65113
rect 263829 65051 264139 65085
rect 263829 65023 263877 65051
rect 263905 65023 263939 65051
rect 263967 65023 264001 65051
rect 264029 65023 264063 65051
rect 264091 65023 264139 65051
rect 263829 64989 264139 65023
rect 263829 64961 263877 64989
rect 263905 64961 263939 64989
rect 263967 64961 264001 64989
rect 264029 64961 264063 64989
rect 264091 64961 264139 64989
rect 263829 56175 264139 64961
rect 263829 56147 263877 56175
rect 263905 56147 263939 56175
rect 263967 56147 264001 56175
rect 264029 56147 264063 56175
rect 264091 56147 264139 56175
rect 263829 56113 264139 56147
rect 263829 56085 263877 56113
rect 263905 56085 263939 56113
rect 263967 56085 264001 56113
rect 264029 56085 264063 56113
rect 264091 56085 264139 56113
rect 263829 56051 264139 56085
rect 263829 56023 263877 56051
rect 263905 56023 263939 56051
rect 263967 56023 264001 56051
rect 264029 56023 264063 56051
rect 264091 56023 264139 56051
rect 263829 55989 264139 56023
rect 263829 55961 263877 55989
rect 263905 55961 263939 55989
rect 263967 55961 264001 55989
rect 264029 55961 264063 55989
rect 264091 55961 264139 55989
rect 263829 47175 264139 55961
rect 263829 47147 263877 47175
rect 263905 47147 263939 47175
rect 263967 47147 264001 47175
rect 264029 47147 264063 47175
rect 264091 47147 264139 47175
rect 263829 47113 264139 47147
rect 263829 47085 263877 47113
rect 263905 47085 263939 47113
rect 263967 47085 264001 47113
rect 264029 47085 264063 47113
rect 264091 47085 264139 47113
rect 263829 47051 264139 47085
rect 263829 47023 263877 47051
rect 263905 47023 263939 47051
rect 263967 47023 264001 47051
rect 264029 47023 264063 47051
rect 264091 47023 264139 47051
rect 263829 46989 264139 47023
rect 263829 46961 263877 46989
rect 263905 46961 263939 46989
rect 263967 46961 264001 46989
rect 264029 46961 264063 46989
rect 264091 46961 264139 46989
rect 263829 38175 264139 46961
rect 263829 38147 263877 38175
rect 263905 38147 263939 38175
rect 263967 38147 264001 38175
rect 264029 38147 264063 38175
rect 264091 38147 264139 38175
rect 263829 38113 264139 38147
rect 263829 38085 263877 38113
rect 263905 38085 263939 38113
rect 263967 38085 264001 38113
rect 264029 38085 264063 38113
rect 264091 38085 264139 38113
rect 263829 38051 264139 38085
rect 263829 38023 263877 38051
rect 263905 38023 263939 38051
rect 263967 38023 264001 38051
rect 264029 38023 264063 38051
rect 264091 38023 264139 38051
rect 263829 37989 264139 38023
rect 263829 37961 263877 37989
rect 263905 37961 263939 37989
rect 263967 37961 264001 37989
rect 264029 37961 264063 37989
rect 264091 37961 264139 37989
rect 263829 29175 264139 37961
rect 263829 29147 263877 29175
rect 263905 29147 263939 29175
rect 263967 29147 264001 29175
rect 264029 29147 264063 29175
rect 264091 29147 264139 29175
rect 263829 29113 264139 29147
rect 263829 29085 263877 29113
rect 263905 29085 263939 29113
rect 263967 29085 264001 29113
rect 264029 29085 264063 29113
rect 264091 29085 264139 29113
rect 263829 29051 264139 29085
rect 263829 29023 263877 29051
rect 263905 29023 263939 29051
rect 263967 29023 264001 29051
rect 264029 29023 264063 29051
rect 264091 29023 264139 29051
rect 263829 28989 264139 29023
rect 263829 28961 263877 28989
rect 263905 28961 263939 28989
rect 263967 28961 264001 28989
rect 264029 28961 264063 28989
rect 264091 28961 264139 28989
rect 263829 20175 264139 28961
rect 263829 20147 263877 20175
rect 263905 20147 263939 20175
rect 263967 20147 264001 20175
rect 264029 20147 264063 20175
rect 264091 20147 264139 20175
rect 263829 20113 264139 20147
rect 263829 20085 263877 20113
rect 263905 20085 263939 20113
rect 263967 20085 264001 20113
rect 264029 20085 264063 20113
rect 264091 20085 264139 20113
rect 263829 20051 264139 20085
rect 263829 20023 263877 20051
rect 263905 20023 263939 20051
rect 263967 20023 264001 20051
rect 264029 20023 264063 20051
rect 264091 20023 264139 20051
rect 263829 19989 264139 20023
rect 263829 19961 263877 19989
rect 263905 19961 263939 19989
rect 263967 19961 264001 19989
rect 264029 19961 264063 19989
rect 264091 19961 264139 19989
rect 263829 11175 264139 19961
rect 263829 11147 263877 11175
rect 263905 11147 263939 11175
rect 263967 11147 264001 11175
rect 264029 11147 264063 11175
rect 264091 11147 264139 11175
rect 263829 11113 264139 11147
rect 263829 11085 263877 11113
rect 263905 11085 263939 11113
rect 263967 11085 264001 11113
rect 264029 11085 264063 11113
rect 264091 11085 264139 11113
rect 263829 11051 264139 11085
rect 263829 11023 263877 11051
rect 263905 11023 263939 11051
rect 263967 11023 264001 11051
rect 264029 11023 264063 11051
rect 264091 11023 264139 11051
rect 263829 10989 264139 11023
rect 263829 10961 263877 10989
rect 263905 10961 263939 10989
rect 263967 10961 264001 10989
rect 264029 10961 264063 10989
rect 264091 10961 264139 10989
rect 263829 2175 264139 10961
rect 263829 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 264139 2175
rect 263829 2113 264139 2147
rect 263829 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 264139 2113
rect 263829 2051 264139 2085
rect 263829 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 264139 2051
rect 263829 1989 264139 2023
rect 263829 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 264139 1989
rect 263829 -80 264139 1961
rect 263829 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 264139 -80
rect 263829 -142 264139 -108
rect 263829 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 264139 -142
rect 263829 -204 264139 -170
rect 263829 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 264139 -204
rect 263829 -266 264139 -232
rect 263829 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 264139 -266
rect 263829 -822 264139 -294
rect 265689 95175 265999 100689
rect 265689 95147 265737 95175
rect 265765 95147 265799 95175
rect 265827 95147 265861 95175
rect 265889 95147 265923 95175
rect 265951 95147 265999 95175
rect 265689 95113 265999 95147
rect 265689 95085 265737 95113
rect 265765 95085 265799 95113
rect 265827 95085 265861 95113
rect 265889 95085 265923 95113
rect 265951 95085 265999 95113
rect 265689 95051 265999 95085
rect 265689 95023 265737 95051
rect 265765 95023 265799 95051
rect 265827 95023 265861 95051
rect 265889 95023 265923 95051
rect 265951 95023 265999 95051
rect 265689 94989 265999 95023
rect 265689 94961 265737 94989
rect 265765 94961 265799 94989
rect 265827 94961 265861 94989
rect 265889 94961 265923 94989
rect 265951 94961 265999 94989
rect 265689 86175 265999 94961
rect 265689 86147 265737 86175
rect 265765 86147 265799 86175
rect 265827 86147 265861 86175
rect 265889 86147 265923 86175
rect 265951 86147 265999 86175
rect 265689 86113 265999 86147
rect 265689 86085 265737 86113
rect 265765 86085 265799 86113
rect 265827 86085 265861 86113
rect 265889 86085 265923 86113
rect 265951 86085 265999 86113
rect 265689 86051 265999 86085
rect 265689 86023 265737 86051
rect 265765 86023 265799 86051
rect 265827 86023 265861 86051
rect 265889 86023 265923 86051
rect 265951 86023 265999 86051
rect 265689 85989 265999 86023
rect 265689 85961 265737 85989
rect 265765 85961 265799 85989
rect 265827 85961 265861 85989
rect 265889 85961 265923 85989
rect 265951 85961 265999 85989
rect 265689 77175 265999 85961
rect 265689 77147 265737 77175
rect 265765 77147 265799 77175
rect 265827 77147 265861 77175
rect 265889 77147 265923 77175
rect 265951 77147 265999 77175
rect 265689 77113 265999 77147
rect 265689 77085 265737 77113
rect 265765 77085 265799 77113
rect 265827 77085 265861 77113
rect 265889 77085 265923 77113
rect 265951 77085 265999 77113
rect 265689 77051 265999 77085
rect 265689 77023 265737 77051
rect 265765 77023 265799 77051
rect 265827 77023 265861 77051
rect 265889 77023 265923 77051
rect 265951 77023 265999 77051
rect 265689 76989 265999 77023
rect 265689 76961 265737 76989
rect 265765 76961 265799 76989
rect 265827 76961 265861 76989
rect 265889 76961 265923 76989
rect 265951 76961 265999 76989
rect 265689 68175 265999 76961
rect 265689 68147 265737 68175
rect 265765 68147 265799 68175
rect 265827 68147 265861 68175
rect 265889 68147 265923 68175
rect 265951 68147 265999 68175
rect 265689 68113 265999 68147
rect 265689 68085 265737 68113
rect 265765 68085 265799 68113
rect 265827 68085 265861 68113
rect 265889 68085 265923 68113
rect 265951 68085 265999 68113
rect 265689 68051 265999 68085
rect 265689 68023 265737 68051
rect 265765 68023 265799 68051
rect 265827 68023 265861 68051
rect 265889 68023 265923 68051
rect 265951 68023 265999 68051
rect 265689 67989 265999 68023
rect 265689 67961 265737 67989
rect 265765 67961 265799 67989
rect 265827 67961 265861 67989
rect 265889 67961 265923 67989
rect 265951 67961 265999 67989
rect 265689 59175 265999 67961
rect 265689 59147 265737 59175
rect 265765 59147 265799 59175
rect 265827 59147 265861 59175
rect 265889 59147 265923 59175
rect 265951 59147 265999 59175
rect 265689 59113 265999 59147
rect 265689 59085 265737 59113
rect 265765 59085 265799 59113
rect 265827 59085 265861 59113
rect 265889 59085 265923 59113
rect 265951 59085 265999 59113
rect 265689 59051 265999 59085
rect 265689 59023 265737 59051
rect 265765 59023 265799 59051
rect 265827 59023 265861 59051
rect 265889 59023 265923 59051
rect 265951 59023 265999 59051
rect 265689 58989 265999 59023
rect 265689 58961 265737 58989
rect 265765 58961 265799 58989
rect 265827 58961 265861 58989
rect 265889 58961 265923 58989
rect 265951 58961 265999 58989
rect 265689 50175 265999 58961
rect 265689 50147 265737 50175
rect 265765 50147 265799 50175
rect 265827 50147 265861 50175
rect 265889 50147 265923 50175
rect 265951 50147 265999 50175
rect 265689 50113 265999 50147
rect 265689 50085 265737 50113
rect 265765 50085 265799 50113
rect 265827 50085 265861 50113
rect 265889 50085 265923 50113
rect 265951 50085 265999 50113
rect 265689 50051 265999 50085
rect 265689 50023 265737 50051
rect 265765 50023 265799 50051
rect 265827 50023 265861 50051
rect 265889 50023 265923 50051
rect 265951 50023 265999 50051
rect 265689 49989 265999 50023
rect 265689 49961 265737 49989
rect 265765 49961 265799 49989
rect 265827 49961 265861 49989
rect 265889 49961 265923 49989
rect 265951 49961 265999 49989
rect 265689 41175 265999 49961
rect 265689 41147 265737 41175
rect 265765 41147 265799 41175
rect 265827 41147 265861 41175
rect 265889 41147 265923 41175
rect 265951 41147 265999 41175
rect 265689 41113 265999 41147
rect 265689 41085 265737 41113
rect 265765 41085 265799 41113
rect 265827 41085 265861 41113
rect 265889 41085 265923 41113
rect 265951 41085 265999 41113
rect 265689 41051 265999 41085
rect 265689 41023 265737 41051
rect 265765 41023 265799 41051
rect 265827 41023 265861 41051
rect 265889 41023 265923 41051
rect 265951 41023 265999 41051
rect 265689 40989 265999 41023
rect 265689 40961 265737 40989
rect 265765 40961 265799 40989
rect 265827 40961 265861 40989
rect 265889 40961 265923 40989
rect 265951 40961 265999 40989
rect 265689 32175 265999 40961
rect 265689 32147 265737 32175
rect 265765 32147 265799 32175
rect 265827 32147 265861 32175
rect 265889 32147 265923 32175
rect 265951 32147 265999 32175
rect 265689 32113 265999 32147
rect 265689 32085 265737 32113
rect 265765 32085 265799 32113
rect 265827 32085 265861 32113
rect 265889 32085 265923 32113
rect 265951 32085 265999 32113
rect 265689 32051 265999 32085
rect 265689 32023 265737 32051
rect 265765 32023 265799 32051
rect 265827 32023 265861 32051
rect 265889 32023 265923 32051
rect 265951 32023 265999 32051
rect 265689 31989 265999 32023
rect 265689 31961 265737 31989
rect 265765 31961 265799 31989
rect 265827 31961 265861 31989
rect 265889 31961 265923 31989
rect 265951 31961 265999 31989
rect 265689 23175 265999 31961
rect 265689 23147 265737 23175
rect 265765 23147 265799 23175
rect 265827 23147 265861 23175
rect 265889 23147 265923 23175
rect 265951 23147 265999 23175
rect 265689 23113 265999 23147
rect 265689 23085 265737 23113
rect 265765 23085 265799 23113
rect 265827 23085 265861 23113
rect 265889 23085 265923 23113
rect 265951 23085 265999 23113
rect 265689 23051 265999 23085
rect 265689 23023 265737 23051
rect 265765 23023 265799 23051
rect 265827 23023 265861 23051
rect 265889 23023 265923 23051
rect 265951 23023 265999 23051
rect 265689 22989 265999 23023
rect 265689 22961 265737 22989
rect 265765 22961 265799 22989
rect 265827 22961 265861 22989
rect 265889 22961 265923 22989
rect 265951 22961 265999 22989
rect 265689 14175 265999 22961
rect 265689 14147 265737 14175
rect 265765 14147 265799 14175
rect 265827 14147 265861 14175
rect 265889 14147 265923 14175
rect 265951 14147 265999 14175
rect 265689 14113 265999 14147
rect 265689 14085 265737 14113
rect 265765 14085 265799 14113
rect 265827 14085 265861 14113
rect 265889 14085 265923 14113
rect 265951 14085 265999 14113
rect 265689 14051 265999 14085
rect 265689 14023 265737 14051
rect 265765 14023 265799 14051
rect 265827 14023 265861 14051
rect 265889 14023 265923 14051
rect 265951 14023 265999 14051
rect 265689 13989 265999 14023
rect 265689 13961 265737 13989
rect 265765 13961 265799 13989
rect 265827 13961 265861 13989
rect 265889 13961 265923 13989
rect 265951 13961 265999 13989
rect 265689 5175 265999 13961
rect 265689 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 265999 5175
rect 265689 5113 265999 5147
rect 265689 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 265999 5113
rect 265689 5051 265999 5085
rect 265689 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 265999 5051
rect 265689 4989 265999 5023
rect 265689 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 265999 4989
rect 265689 -560 265999 4961
rect 265689 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 265999 -560
rect 265689 -622 265999 -588
rect 265689 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 265999 -622
rect 265689 -684 265999 -650
rect 265689 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 265999 -684
rect 265689 -746 265999 -712
rect 265689 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 265999 -746
rect 265689 -822 265999 -774
rect 279189 92175 279499 100961
rect 279189 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 279499 92175
rect 279189 92113 279499 92147
rect 279189 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 279499 92113
rect 279189 92051 279499 92085
rect 279189 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 279499 92051
rect 279189 91989 279499 92023
rect 279189 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 279499 91989
rect 279189 83175 279499 91961
rect 279189 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 279499 83175
rect 279189 83113 279499 83147
rect 279189 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 279499 83113
rect 279189 83051 279499 83085
rect 279189 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 279499 83051
rect 279189 82989 279499 83023
rect 279189 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 279499 82989
rect 279189 74175 279499 82961
rect 279189 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 279499 74175
rect 279189 74113 279499 74147
rect 279189 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 279499 74113
rect 279189 74051 279499 74085
rect 279189 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 279499 74051
rect 279189 73989 279499 74023
rect 279189 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 279499 73989
rect 279189 65175 279499 73961
rect 279189 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 279499 65175
rect 279189 65113 279499 65147
rect 279189 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 279499 65113
rect 279189 65051 279499 65085
rect 279189 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 279499 65051
rect 279189 64989 279499 65023
rect 279189 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 279499 64989
rect 279189 56175 279499 64961
rect 279189 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 279499 56175
rect 279189 56113 279499 56147
rect 279189 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 279499 56113
rect 279189 56051 279499 56085
rect 279189 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 279499 56051
rect 279189 55989 279499 56023
rect 279189 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 279499 55989
rect 279189 47175 279499 55961
rect 279189 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 279499 47175
rect 279189 47113 279499 47147
rect 279189 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 279499 47113
rect 279189 47051 279499 47085
rect 279189 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 279499 47051
rect 279189 46989 279499 47023
rect 279189 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 279499 46989
rect 279189 38175 279499 46961
rect 279189 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 279499 38175
rect 279189 38113 279499 38147
rect 279189 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 279499 38113
rect 279189 38051 279499 38085
rect 279189 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 279499 38051
rect 279189 37989 279499 38023
rect 279189 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 279499 37989
rect 279189 29175 279499 37961
rect 279189 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 279499 29175
rect 279189 29113 279499 29147
rect 279189 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 279499 29113
rect 279189 29051 279499 29085
rect 279189 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 279499 29051
rect 279189 28989 279499 29023
rect 279189 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 279499 28989
rect 279189 20175 279499 28961
rect 279189 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 279499 20175
rect 279189 20113 279499 20147
rect 279189 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 279499 20113
rect 279189 20051 279499 20085
rect 279189 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 279499 20051
rect 279189 19989 279499 20023
rect 279189 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 279499 19989
rect 279189 11175 279499 19961
rect 279189 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 279499 11175
rect 279189 11113 279499 11147
rect 279189 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 279499 11113
rect 279189 11051 279499 11085
rect 279189 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 279499 11051
rect 279189 10989 279499 11023
rect 279189 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 279499 10989
rect 279189 2175 279499 10961
rect 279189 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 279499 2175
rect 279189 2113 279499 2147
rect 279189 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 279499 2113
rect 279189 2051 279499 2085
rect 279189 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 279499 2051
rect 279189 1989 279499 2023
rect 279189 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 279499 1989
rect 279189 -80 279499 1961
rect 279189 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 279499 -80
rect 279189 -142 279499 -108
rect 279189 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 279499 -142
rect 279189 -204 279499 -170
rect 279189 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 279499 -204
rect 279189 -266 279499 -232
rect 279189 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 279499 -266
rect 279189 -822 279499 -294
rect 281049 299086 281359 299134
rect 281049 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 281359 299086
rect 281049 299024 281359 299058
rect 281049 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 281359 299024
rect 281049 298962 281359 298996
rect 281049 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 281359 298962
rect 281049 298900 281359 298934
rect 281049 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 281359 298900
rect 281049 293175 281359 298872
rect 281049 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 281359 293175
rect 281049 293113 281359 293147
rect 281049 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 281359 293113
rect 281049 293051 281359 293085
rect 281049 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 281359 293051
rect 281049 292989 281359 293023
rect 281049 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 281359 292989
rect 281049 284175 281359 292961
rect 281049 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 281359 284175
rect 281049 284113 281359 284147
rect 281049 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 281359 284113
rect 281049 284051 281359 284085
rect 281049 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 281359 284051
rect 281049 283989 281359 284023
rect 281049 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 281359 283989
rect 281049 275175 281359 283961
rect 281049 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 281359 275175
rect 281049 275113 281359 275147
rect 281049 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 281359 275113
rect 281049 275051 281359 275085
rect 281049 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 281359 275051
rect 281049 274989 281359 275023
rect 294549 298606 294859 299134
rect 294549 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 294859 298606
rect 294549 298544 294859 298578
rect 294549 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 294859 298544
rect 294549 298482 294859 298516
rect 294549 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 294859 298482
rect 294549 298420 294859 298454
rect 294549 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 294859 298420
rect 294549 290175 294859 298392
rect 294549 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 294859 290175
rect 294549 290113 294859 290147
rect 294549 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 294859 290113
rect 294549 290051 294859 290085
rect 294549 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 294859 290051
rect 294549 289989 294859 290023
rect 294549 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 294859 289989
rect 294549 281175 294859 289961
rect 294549 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 294859 281175
rect 294549 281113 294859 281147
rect 294549 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 294859 281113
rect 294549 281051 294859 281085
rect 294549 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 294859 281051
rect 294549 280989 294859 281023
rect 294549 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 294859 280989
rect 281049 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 281359 274989
rect 281049 266175 281359 274961
rect 281049 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 281359 266175
rect 281049 266113 281359 266147
rect 281049 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 281359 266113
rect 281049 266051 281359 266085
rect 281049 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 281359 266051
rect 281049 265989 281359 266023
rect 281049 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 281359 265989
rect 281049 257175 281359 265961
rect 281049 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 281359 257175
rect 281049 257113 281359 257147
rect 281049 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 281359 257113
rect 281049 257051 281359 257085
rect 281049 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 281359 257051
rect 281049 256989 281359 257023
rect 281049 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 281359 256989
rect 281049 248175 281359 256961
rect 281049 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 281359 248175
rect 281049 248113 281359 248147
rect 281049 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 281359 248113
rect 281049 248051 281359 248085
rect 281049 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 281359 248051
rect 281049 247989 281359 248023
rect 281049 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 281359 247989
rect 281049 239175 281359 247961
rect 281049 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 281359 239175
rect 281049 239113 281359 239147
rect 281049 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 281359 239113
rect 281049 239051 281359 239085
rect 281049 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 281359 239051
rect 281049 238989 281359 239023
rect 281049 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 281359 238989
rect 281049 230175 281359 238961
rect 281049 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 281359 230175
rect 281049 230113 281359 230147
rect 281049 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 281359 230113
rect 281049 230051 281359 230085
rect 281049 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 281359 230051
rect 281049 229989 281359 230023
rect 281049 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 281359 229989
rect 281049 221175 281359 229961
rect 281049 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 281359 221175
rect 281049 221113 281359 221147
rect 281049 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 281359 221113
rect 281049 221051 281359 221085
rect 281049 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 281359 221051
rect 281049 220989 281359 221023
rect 281049 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 281359 220989
rect 281049 212175 281359 220961
rect 281049 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 281359 212175
rect 281049 212113 281359 212147
rect 281049 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 281359 212113
rect 281049 212051 281359 212085
rect 281049 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 281359 212051
rect 281049 211989 281359 212023
rect 281049 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 281359 211989
rect 281049 203175 281359 211961
rect 281049 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 281359 203175
rect 281049 203113 281359 203147
rect 281049 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 281359 203113
rect 281049 203051 281359 203085
rect 281049 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 281359 203051
rect 281049 202989 281359 203023
rect 281049 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 281359 202989
rect 281049 194175 281359 202961
rect 281049 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 281359 194175
rect 281049 194113 281359 194147
rect 281049 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 281359 194113
rect 281049 194051 281359 194085
rect 281049 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 281359 194051
rect 281049 193989 281359 194023
rect 281049 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 281359 193989
rect 281049 185175 281359 193961
rect 281049 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 281359 185175
rect 281049 185113 281359 185147
rect 281049 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 281359 185113
rect 281049 185051 281359 185085
rect 281049 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 281359 185051
rect 281049 184989 281359 185023
rect 281049 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 281359 184989
rect 281049 176175 281359 184961
rect 281049 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 281359 176175
rect 281049 176113 281359 176147
rect 281049 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 281359 176113
rect 281049 176051 281359 176085
rect 281049 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 281359 176051
rect 281049 175989 281359 176023
rect 281049 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 281359 175989
rect 281049 167175 281359 175961
rect 281049 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 281359 167175
rect 281049 167113 281359 167147
rect 281049 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 281359 167113
rect 281049 167051 281359 167085
rect 281049 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 281359 167051
rect 281049 166989 281359 167023
rect 281049 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 281359 166989
rect 281049 158175 281359 166961
rect 281049 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 281359 158175
rect 281049 158113 281359 158147
rect 281049 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 281359 158113
rect 281049 158051 281359 158085
rect 281049 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 281359 158051
rect 281049 157989 281359 158023
rect 281049 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 281359 157989
rect 281049 149175 281359 157961
rect 281414 275002 281442 275007
rect 281414 156338 281442 274974
rect 294549 272175 294859 280961
rect 294549 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 294859 272175
rect 294549 272113 294859 272147
rect 294549 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 294859 272113
rect 294549 272051 294859 272085
rect 294549 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 294859 272051
rect 294549 271989 294859 272023
rect 294549 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 294859 271989
rect 281806 267610 281834 267615
rect 281414 156305 281442 156310
rect 281470 238042 281498 238047
rect 281049 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 281359 149175
rect 281049 149113 281359 149147
rect 281049 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 281359 149113
rect 281049 149051 281359 149085
rect 281049 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 281359 149051
rect 281049 148989 281359 149023
rect 281049 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 281359 148989
rect 281049 140175 281359 148961
rect 281049 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 281359 140175
rect 281049 140113 281359 140147
rect 281049 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 281359 140113
rect 281049 140051 281359 140085
rect 281049 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 281359 140051
rect 281049 139989 281359 140023
rect 281049 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 281359 139989
rect 281049 131175 281359 139961
rect 281049 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 281359 131175
rect 281049 131113 281359 131147
rect 281049 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 281359 131113
rect 281049 131051 281359 131085
rect 281049 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 281359 131051
rect 281049 130989 281359 131023
rect 281049 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 281359 130989
rect 281049 122175 281359 130961
rect 281470 126882 281498 238014
rect 281470 126849 281498 126854
rect 281526 215866 281554 215871
rect 281049 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 281359 122175
rect 281049 122113 281359 122147
rect 281049 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 281359 122113
rect 281049 122051 281359 122085
rect 281049 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 281359 122051
rect 281049 121989 281359 122023
rect 281049 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 281359 121989
rect 281049 113175 281359 121961
rect 281526 119322 281554 215838
rect 281526 119289 281554 119294
rect 281582 193690 281610 193695
rect 281049 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 281359 113175
rect 281049 113113 281359 113147
rect 281049 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 281359 113113
rect 281049 113051 281359 113085
rect 281049 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 281359 113051
rect 281049 112989 281359 113023
rect 281049 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 281359 112989
rect 281049 104175 281359 112961
rect 281582 104930 281610 193662
rect 281806 148946 281834 267582
rect 294549 263175 294859 271961
rect 294549 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 294859 263175
rect 294549 263113 294859 263147
rect 294549 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 294859 263113
rect 294549 263051 294859 263085
rect 294549 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 294859 263051
rect 294549 262989 294859 263023
rect 294549 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 294859 262989
rect 281806 148913 281834 148918
rect 281862 260218 281890 260223
rect 281862 142338 281890 260190
rect 294549 254175 294859 262961
rect 294549 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 294859 254175
rect 294549 254113 294859 254147
rect 294549 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 294859 254113
rect 294549 254051 294859 254085
rect 294549 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 294859 254051
rect 294549 253989 294859 254023
rect 294549 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 294859 253989
rect 284326 252826 284354 252831
rect 283486 230650 283514 230655
rect 282646 208474 282674 208479
rect 281862 142305 281890 142310
rect 281918 186298 281946 186303
rect 281806 141946 281834 141951
rect 281582 104897 281610 104902
rect 281750 104986 281778 104991
rect 281049 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 281359 104175
rect 281049 104113 281359 104147
rect 281049 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 281359 104113
rect 281049 104051 281359 104085
rect 281049 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 281359 104051
rect 281049 103989 281359 104023
rect 281049 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 281359 103989
rect 281049 95175 281359 103961
rect 281049 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 281359 95175
rect 281049 95113 281359 95147
rect 281049 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 281359 95113
rect 281049 95051 281359 95085
rect 281049 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 281359 95051
rect 281049 94989 281359 95023
rect 281049 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 281359 94989
rect 281049 86175 281359 94961
rect 281049 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 281359 86175
rect 281049 86113 281359 86147
rect 281049 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 281359 86113
rect 281049 86051 281359 86085
rect 281049 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 281359 86051
rect 281049 85989 281359 86023
rect 281049 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 281359 85989
rect 281049 77175 281359 85961
rect 281049 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 281359 77175
rect 281049 77113 281359 77147
rect 281049 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 281359 77113
rect 281049 77051 281359 77085
rect 281049 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 281359 77051
rect 281049 76989 281359 77023
rect 281049 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 281359 76989
rect 281049 68175 281359 76961
rect 281049 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 281359 68175
rect 281049 68113 281359 68147
rect 281049 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 281359 68113
rect 281049 68051 281359 68085
rect 281049 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 281359 68051
rect 281049 67989 281359 68023
rect 281049 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 281359 67989
rect 281049 59175 281359 67961
rect 281049 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 281359 59175
rect 281049 59113 281359 59147
rect 281049 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 281359 59113
rect 281049 59051 281359 59085
rect 281049 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 281359 59051
rect 281049 58989 281359 59023
rect 281049 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 281359 58989
rect 281049 50175 281359 58961
rect 281049 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 281359 50175
rect 281049 50113 281359 50147
rect 281049 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 281359 50113
rect 281049 50051 281359 50085
rect 281049 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 281359 50051
rect 281049 49989 281359 50023
rect 281049 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 281359 49989
rect 281049 41175 281359 49961
rect 281049 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 281359 41175
rect 281049 41113 281359 41147
rect 281049 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 281359 41113
rect 281049 41051 281359 41085
rect 281049 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 281359 41051
rect 281049 40989 281359 41023
rect 281049 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 281359 40989
rect 281049 32175 281359 40961
rect 281049 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 281359 32175
rect 281049 32113 281359 32147
rect 281049 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 281359 32113
rect 281049 32051 281359 32085
rect 281049 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 281359 32051
rect 281049 31989 281359 32023
rect 281049 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 281359 31989
rect 281049 23175 281359 31961
rect 281049 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 281359 23175
rect 281049 23113 281359 23147
rect 281049 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 281359 23113
rect 281049 23051 281359 23085
rect 281049 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 281359 23051
rect 281049 22989 281359 23023
rect 281049 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 281359 22989
rect 281049 14175 281359 22961
rect 281049 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 281359 14175
rect 281049 14113 281359 14147
rect 281049 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 281359 14113
rect 281049 14051 281359 14085
rect 281049 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 281359 14051
rect 281049 13989 281359 14023
rect 281049 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 281359 13989
rect 281049 5175 281359 13961
rect 281049 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 281359 5175
rect 281049 5113 281359 5147
rect 281049 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 281359 5113
rect 281049 5051 281359 5085
rect 281049 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 281359 5051
rect 281049 4989 281359 5023
rect 281049 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 281359 4989
rect 281049 -560 281359 4961
rect 281750 3570 281778 104958
rect 281806 36610 281834 141918
rect 281806 36577 281834 36582
rect 281862 127162 281890 127167
rect 281862 23394 281890 127134
rect 281918 76258 281946 186270
rect 281918 76225 281946 76230
rect 281974 171514 282002 171519
rect 281974 63042 282002 171486
rect 281974 63009 282002 63014
rect 282030 164122 282058 164127
rect 282030 56434 282058 164094
rect 282030 56401 282058 56406
rect 282086 156730 282114 156735
rect 282086 49826 282114 156702
rect 282086 49793 282114 49798
rect 282142 149338 282170 149343
rect 282142 43218 282170 149310
rect 282142 43185 282170 43190
rect 282198 119770 282226 119775
rect 281862 23361 281890 23366
rect 282198 16842 282226 119742
rect 282646 96082 282674 208446
rect 283486 115962 283514 230622
rect 284326 135730 284354 252798
rect 286846 245434 286874 245439
rect 284326 135697 284354 135702
rect 286006 223258 286034 223263
rect 283486 115929 283514 115934
rect 282646 96049 282674 96054
rect 285166 112378 285194 112383
rect 282198 16809 282226 16814
rect 285166 10178 285194 112350
rect 286006 109298 286034 223230
rect 286846 129122 286874 245406
rect 294549 245175 294859 253961
rect 294549 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 294859 245175
rect 294549 245113 294859 245147
rect 294549 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 294859 245113
rect 294549 245051 294859 245085
rect 294549 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 294859 245051
rect 294549 244989 294859 245023
rect 294549 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 294859 244989
rect 294549 236175 294859 244961
rect 294549 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 294859 236175
rect 294549 236113 294859 236147
rect 294549 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 294859 236113
rect 294549 236051 294859 236085
rect 294549 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 294859 236051
rect 294549 235989 294859 236023
rect 294549 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 294859 235989
rect 294549 227175 294859 235961
rect 294549 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 294859 227175
rect 294549 227113 294859 227147
rect 294549 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 294859 227113
rect 294549 227051 294859 227085
rect 294549 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 294859 227051
rect 294549 226989 294859 227023
rect 294549 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 294859 226989
rect 294549 218175 294859 226961
rect 294549 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 294859 218175
rect 294549 218113 294859 218147
rect 294549 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 294859 218113
rect 294549 218051 294859 218085
rect 294549 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 294859 218051
rect 294549 217989 294859 218023
rect 294549 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 294859 217989
rect 294549 209175 294859 217961
rect 294549 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 294859 209175
rect 294549 209113 294859 209147
rect 294549 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 294859 209113
rect 294549 209051 294859 209085
rect 294549 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 294859 209051
rect 294549 208989 294859 209023
rect 294549 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 294859 208989
rect 292726 201082 292754 201087
rect 289366 178906 289394 178911
rect 286846 129089 286874 129094
rect 287686 134554 287714 134559
rect 286006 109265 286034 109270
rect 287686 30002 287714 134526
rect 289366 69650 289394 178878
rect 292726 89586 292754 201054
rect 292726 89553 292754 89558
rect 294549 200175 294859 208961
rect 294549 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 294859 200175
rect 294549 200113 294859 200147
rect 294549 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 294859 200113
rect 294549 200051 294859 200085
rect 294549 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 294859 200051
rect 294549 199989 294859 200023
rect 294549 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 294859 199989
rect 294549 191175 294859 199961
rect 294549 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 294859 191175
rect 294549 191113 294859 191147
rect 294549 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 294859 191113
rect 294549 191051 294859 191085
rect 294549 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 294859 191051
rect 294549 190989 294859 191023
rect 294549 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 294859 190989
rect 294549 182175 294859 190961
rect 294549 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 294859 182175
rect 294549 182113 294859 182147
rect 294549 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 294859 182113
rect 294549 182051 294859 182085
rect 294549 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 294859 182051
rect 294549 181989 294859 182023
rect 294549 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 294859 181989
rect 294549 173175 294859 181961
rect 294549 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 294859 173175
rect 294549 173113 294859 173147
rect 294549 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 294859 173113
rect 294549 173051 294859 173085
rect 294549 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 294859 173051
rect 294549 172989 294859 173023
rect 294549 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 294859 172989
rect 294549 164175 294859 172961
rect 294549 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 294859 164175
rect 294549 164113 294859 164147
rect 294549 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 294859 164113
rect 294549 164051 294859 164085
rect 294549 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 294859 164051
rect 294549 163989 294859 164023
rect 294549 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 294859 163989
rect 294549 155175 294859 163961
rect 294549 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 294859 155175
rect 294549 155113 294859 155147
rect 294549 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 294859 155113
rect 294549 155051 294859 155085
rect 294549 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 294859 155051
rect 294549 154989 294859 155023
rect 294549 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 294859 154989
rect 294549 146175 294859 154961
rect 294549 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 294859 146175
rect 294549 146113 294859 146147
rect 294549 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 294859 146113
rect 294549 146051 294859 146085
rect 294549 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 294859 146051
rect 294549 145989 294859 146023
rect 294549 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 294859 145989
rect 294549 137175 294859 145961
rect 294549 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 294859 137175
rect 294549 137113 294859 137147
rect 294549 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 294859 137113
rect 294549 137051 294859 137085
rect 294549 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 294859 137051
rect 294549 136989 294859 137023
rect 294549 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 294859 136989
rect 294549 128175 294859 136961
rect 294549 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 294859 128175
rect 294549 128113 294859 128147
rect 294549 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 294859 128113
rect 294549 128051 294859 128085
rect 294549 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 294859 128051
rect 294549 127989 294859 128023
rect 294549 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 294859 127989
rect 294549 119175 294859 127961
rect 294549 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 294859 119175
rect 294549 119113 294859 119147
rect 294549 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 294859 119113
rect 294549 119051 294859 119085
rect 294549 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 294859 119051
rect 294549 118989 294859 119023
rect 294549 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 294859 118989
rect 294549 110175 294859 118961
rect 294549 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 294859 110175
rect 294549 110113 294859 110147
rect 294549 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 294859 110113
rect 294549 110051 294859 110085
rect 294549 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 294859 110051
rect 294549 109989 294859 110023
rect 294549 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 294859 109989
rect 294549 101175 294859 109961
rect 294549 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 294859 101175
rect 294549 101113 294859 101147
rect 294549 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 294859 101113
rect 294549 101051 294859 101085
rect 294549 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 294859 101051
rect 294549 100989 294859 101023
rect 294549 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 294859 100989
rect 294549 92175 294859 100961
rect 294549 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 294859 92175
rect 294549 92113 294859 92147
rect 294549 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 294859 92113
rect 294549 92051 294859 92085
rect 294549 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 294859 92051
rect 294549 91989 294859 92023
rect 294549 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 294859 91989
rect 289366 69617 289394 69622
rect 294549 83175 294859 91961
rect 294549 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 294859 83175
rect 294549 83113 294859 83147
rect 294549 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 294859 83113
rect 294549 83051 294859 83085
rect 294549 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 294859 83051
rect 294549 82989 294859 83023
rect 294549 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 294859 82989
rect 294549 74175 294859 82961
rect 294549 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 294859 74175
rect 294549 74113 294859 74147
rect 294549 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 294859 74113
rect 294549 74051 294859 74085
rect 294549 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 294859 74051
rect 294549 73989 294859 74023
rect 294549 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 294859 73989
rect 287686 29969 287714 29974
rect 294549 65175 294859 73961
rect 294549 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 294859 65175
rect 294549 65113 294859 65147
rect 294549 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 294859 65113
rect 294549 65051 294859 65085
rect 294549 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 294859 65051
rect 294549 64989 294859 65023
rect 294549 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 294859 64989
rect 294549 56175 294859 64961
rect 294549 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 294859 56175
rect 294549 56113 294859 56147
rect 294549 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 294859 56113
rect 294549 56051 294859 56085
rect 294549 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 294859 56051
rect 294549 55989 294859 56023
rect 294549 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 294859 55989
rect 294549 47175 294859 55961
rect 294549 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 294859 47175
rect 294549 47113 294859 47147
rect 294549 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 294859 47113
rect 294549 47051 294859 47085
rect 294549 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 294859 47051
rect 294549 46989 294859 47023
rect 294549 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 294859 46989
rect 294549 38175 294859 46961
rect 294549 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 294859 38175
rect 294549 38113 294859 38147
rect 294549 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 294859 38113
rect 294549 38051 294859 38085
rect 294549 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 294859 38051
rect 294549 37989 294859 38023
rect 294549 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 294859 37989
rect 285166 10145 285194 10150
rect 294549 29175 294859 37961
rect 294549 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 294859 29175
rect 294549 29113 294859 29147
rect 294549 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 294859 29113
rect 294549 29051 294859 29085
rect 294549 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 294859 29051
rect 294549 28989 294859 29023
rect 294549 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 294859 28989
rect 294549 20175 294859 28961
rect 294549 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 294859 20175
rect 294549 20113 294859 20147
rect 294549 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 294859 20113
rect 294549 20051 294859 20085
rect 294549 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 294859 20051
rect 294549 19989 294859 20023
rect 294549 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 294859 19989
rect 294549 11175 294859 19961
rect 294549 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 294859 11175
rect 294549 11113 294859 11147
rect 294549 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 294859 11113
rect 294549 11051 294859 11085
rect 294549 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 294859 11051
rect 294549 10989 294859 11023
rect 294549 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 294859 10989
rect 281750 3537 281778 3542
rect 281049 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 281359 -560
rect 281049 -622 281359 -588
rect 281049 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 281359 -622
rect 281049 -684 281359 -650
rect 281049 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 281359 -684
rect 281049 -746 281359 -712
rect 281049 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 281359 -746
rect 281049 -822 281359 -774
rect 294549 2175 294859 10961
rect 294549 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 294859 2175
rect 294549 2113 294859 2147
rect 294549 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 294859 2113
rect 294549 2051 294859 2085
rect 294549 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 294859 2051
rect 294549 1989 294859 2023
rect 294549 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 294859 1989
rect 294549 -80 294859 1961
rect 294549 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 294859 -80
rect 294549 -142 294859 -108
rect 294549 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 294859 -142
rect 294549 -204 294859 -170
rect 294549 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 294859 -204
rect 294549 -266 294859 -232
rect 294549 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 294859 -266
rect 294549 -822 294859 -294
rect 296409 299086 296719 299134
rect 296409 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 296719 299086
rect 296409 299024 296719 299058
rect 296409 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 296719 299024
rect 296409 298962 296719 298996
rect 296409 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 296719 298962
rect 296409 298900 296719 298934
rect 296409 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 296719 298900
rect 296409 293175 296719 298872
rect 298680 299086 298990 299134
rect 298680 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect 298680 299024 298990 299058
rect 298680 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect 298680 298962 298990 298996
rect 298680 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect 298680 298900 298990 298934
rect 298680 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect 296409 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 296719 293175
rect 296409 293113 296719 293147
rect 296409 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 296719 293113
rect 296409 293051 296719 293085
rect 296409 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 296719 293051
rect 296409 292989 296719 293023
rect 296409 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 296719 292989
rect 296409 284175 296719 292961
rect 296409 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 296719 284175
rect 296409 284113 296719 284147
rect 296409 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 296719 284113
rect 296409 284051 296719 284085
rect 296409 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 296719 284051
rect 296409 283989 296719 284023
rect 296409 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 296719 283989
rect 296409 275175 296719 283961
rect 296409 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 296719 275175
rect 296409 275113 296719 275147
rect 296409 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 296719 275113
rect 296409 275051 296719 275085
rect 296409 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 296719 275051
rect 296409 274989 296719 275023
rect 296409 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 296719 274989
rect 296409 266175 296719 274961
rect 296409 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 296719 266175
rect 296409 266113 296719 266147
rect 296409 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 296719 266113
rect 296409 266051 296719 266085
rect 296409 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 296719 266051
rect 296409 265989 296719 266023
rect 296409 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 296719 265989
rect 296409 257175 296719 265961
rect 296409 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 296719 257175
rect 296409 257113 296719 257147
rect 296409 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 296719 257113
rect 296409 257051 296719 257085
rect 296409 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 296719 257051
rect 296409 256989 296719 257023
rect 296409 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 296719 256989
rect 296409 248175 296719 256961
rect 296409 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 296719 248175
rect 296409 248113 296719 248147
rect 296409 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 296719 248113
rect 296409 248051 296719 248085
rect 296409 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 296719 248051
rect 296409 247989 296719 248023
rect 296409 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 296719 247989
rect 296409 239175 296719 247961
rect 296409 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 296719 239175
rect 296409 239113 296719 239147
rect 296409 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 296719 239113
rect 296409 239051 296719 239085
rect 296409 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 296719 239051
rect 296409 238989 296719 239023
rect 296409 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 296719 238989
rect 296409 230175 296719 238961
rect 296409 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 296719 230175
rect 296409 230113 296719 230147
rect 296409 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 296719 230113
rect 296409 230051 296719 230085
rect 296409 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 296719 230051
rect 296409 229989 296719 230023
rect 296409 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 296719 229989
rect 296409 221175 296719 229961
rect 296409 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 296719 221175
rect 296409 221113 296719 221147
rect 296409 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 296719 221113
rect 296409 221051 296719 221085
rect 296409 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 296719 221051
rect 296409 220989 296719 221023
rect 296409 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 296719 220989
rect 296409 212175 296719 220961
rect 296409 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 296719 212175
rect 296409 212113 296719 212147
rect 296409 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 296719 212113
rect 296409 212051 296719 212085
rect 296409 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 296719 212051
rect 296409 211989 296719 212023
rect 296409 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 296719 211989
rect 296409 203175 296719 211961
rect 296409 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 296719 203175
rect 296409 203113 296719 203147
rect 296409 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 296719 203113
rect 296409 203051 296719 203085
rect 296409 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 296719 203051
rect 296409 202989 296719 203023
rect 296409 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 296719 202989
rect 296409 194175 296719 202961
rect 296409 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 296719 194175
rect 296409 194113 296719 194147
rect 296409 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 296719 194113
rect 296409 194051 296719 194085
rect 296409 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 296719 194051
rect 296409 193989 296719 194023
rect 296409 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 296719 193989
rect 296409 185175 296719 193961
rect 296409 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 296719 185175
rect 296409 185113 296719 185147
rect 296409 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 296719 185113
rect 296409 185051 296719 185085
rect 296409 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 296719 185051
rect 296409 184989 296719 185023
rect 296409 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 296719 184989
rect 296409 176175 296719 184961
rect 296409 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 296719 176175
rect 296409 176113 296719 176147
rect 296409 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 296719 176113
rect 296409 176051 296719 176085
rect 296409 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 296719 176051
rect 296409 175989 296719 176023
rect 296409 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 296719 175989
rect 296409 167175 296719 175961
rect 296409 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 296719 167175
rect 296409 167113 296719 167147
rect 296409 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 296719 167113
rect 296409 167051 296719 167085
rect 296409 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 296719 167051
rect 296409 166989 296719 167023
rect 296409 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 296719 166989
rect 296409 158175 296719 166961
rect 296409 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 296719 158175
rect 296409 158113 296719 158147
rect 296409 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 296719 158113
rect 296409 158051 296719 158085
rect 296409 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 296719 158051
rect 296409 157989 296719 158023
rect 296409 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 296719 157989
rect 296409 149175 296719 157961
rect 296409 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 296719 149175
rect 296409 149113 296719 149147
rect 296409 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 296719 149113
rect 296409 149051 296719 149085
rect 296409 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 296719 149051
rect 296409 148989 296719 149023
rect 296409 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 296719 148989
rect 296409 140175 296719 148961
rect 296409 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 296719 140175
rect 296409 140113 296719 140147
rect 296409 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 296719 140113
rect 296409 140051 296719 140085
rect 296409 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 296719 140051
rect 296409 139989 296719 140023
rect 296409 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 296719 139989
rect 296409 131175 296719 139961
rect 296409 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 296719 131175
rect 296409 131113 296719 131147
rect 296409 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 296719 131113
rect 296409 131051 296719 131085
rect 296409 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 296719 131051
rect 296409 130989 296719 131023
rect 296409 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 296719 130989
rect 296409 122175 296719 130961
rect 296409 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 296719 122175
rect 296409 122113 296719 122147
rect 296409 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 296719 122113
rect 296409 122051 296719 122085
rect 296409 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 296719 122051
rect 296409 121989 296719 122023
rect 296409 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 296719 121989
rect 296409 113175 296719 121961
rect 296409 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 296719 113175
rect 296409 113113 296719 113147
rect 296409 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 296719 113113
rect 296409 113051 296719 113085
rect 296409 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 296719 113051
rect 296409 112989 296719 113023
rect 296409 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 296719 112989
rect 296409 104175 296719 112961
rect 296409 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 296719 104175
rect 296409 104113 296719 104147
rect 296409 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 296719 104113
rect 296409 104051 296719 104085
rect 296409 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 296719 104051
rect 296409 103989 296719 104023
rect 296409 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 296719 103989
rect 296409 95175 296719 103961
rect 296409 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 296719 95175
rect 296409 95113 296719 95147
rect 296409 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 296719 95113
rect 296409 95051 296719 95085
rect 296409 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 296719 95051
rect 296409 94989 296719 95023
rect 296409 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 296719 94989
rect 296409 86175 296719 94961
rect 296409 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 296719 86175
rect 296409 86113 296719 86147
rect 296409 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 296719 86113
rect 296409 86051 296719 86085
rect 296409 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 296719 86051
rect 296409 85989 296719 86023
rect 296409 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 296719 85989
rect 296409 77175 296719 85961
rect 296409 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 296719 77175
rect 296409 77113 296719 77147
rect 296409 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 296719 77113
rect 296409 77051 296719 77085
rect 296409 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 296719 77051
rect 296409 76989 296719 77023
rect 296409 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 296719 76989
rect 296409 68175 296719 76961
rect 296409 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 296719 68175
rect 296409 68113 296719 68147
rect 296409 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 296719 68113
rect 296409 68051 296719 68085
rect 296409 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 296719 68051
rect 296409 67989 296719 68023
rect 296409 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 296719 67989
rect 296409 59175 296719 67961
rect 296409 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 296719 59175
rect 296409 59113 296719 59147
rect 296409 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 296719 59113
rect 296409 59051 296719 59085
rect 296409 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 296719 59051
rect 296409 58989 296719 59023
rect 296409 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 296719 58989
rect 296409 50175 296719 58961
rect 296409 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 296719 50175
rect 296409 50113 296719 50147
rect 296409 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 296719 50113
rect 296409 50051 296719 50085
rect 296409 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 296719 50051
rect 296409 49989 296719 50023
rect 296409 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 296719 49989
rect 296409 41175 296719 49961
rect 296409 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 296719 41175
rect 296409 41113 296719 41147
rect 296409 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 296719 41113
rect 296409 41051 296719 41085
rect 296409 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 296719 41051
rect 296409 40989 296719 41023
rect 296409 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 296719 40989
rect 296409 32175 296719 40961
rect 296409 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 296719 32175
rect 296409 32113 296719 32147
rect 296409 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 296719 32113
rect 296409 32051 296719 32085
rect 296409 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 296719 32051
rect 296409 31989 296719 32023
rect 296409 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 296719 31989
rect 296409 23175 296719 31961
rect 296409 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 296719 23175
rect 296409 23113 296719 23147
rect 296409 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 296719 23113
rect 296409 23051 296719 23085
rect 296409 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 296719 23051
rect 296409 22989 296719 23023
rect 296409 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 296719 22989
rect 296409 14175 296719 22961
rect 296409 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 296719 14175
rect 296409 14113 296719 14147
rect 296409 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 296719 14113
rect 296409 14051 296719 14085
rect 296409 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 296719 14051
rect 296409 13989 296719 14023
rect 296409 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 296719 13989
rect 296409 5175 296719 13961
rect 296409 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 296719 5175
rect 296409 5113 296719 5147
rect 296409 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 296719 5113
rect 296409 5051 296719 5085
rect 296409 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 296719 5051
rect 296409 4989 296719 5023
rect 296409 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 296719 4989
rect 296409 -560 296719 4961
rect 298200 298606 298510 298654
rect 298200 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect 298200 298544 298510 298578
rect 298200 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect 298200 298482 298510 298516
rect 298200 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect 298200 298420 298510 298454
rect 298200 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect 298200 290175 298510 298392
rect 298200 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298510 290175
rect 298200 290113 298510 290147
rect 298200 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298510 290113
rect 298200 290051 298510 290085
rect 298200 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298510 290051
rect 298200 289989 298510 290023
rect 298200 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298510 289989
rect 298200 281175 298510 289961
rect 298200 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298510 281175
rect 298200 281113 298510 281147
rect 298200 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298510 281113
rect 298200 281051 298510 281085
rect 298200 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298510 281051
rect 298200 280989 298510 281023
rect 298200 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298510 280989
rect 298200 272175 298510 280961
rect 298200 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298510 272175
rect 298200 272113 298510 272147
rect 298200 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298510 272113
rect 298200 272051 298510 272085
rect 298200 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298510 272051
rect 298200 271989 298510 272023
rect 298200 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298510 271989
rect 298200 263175 298510 271961
rect 298200 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298510 263175
rect 298200 263113 298510 263147
rect 298200 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298510 263113
rect 298200 263051 298510 263085
rect 298200 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298510 263051
rect 298200 262989 298510 263023
rect 298200 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298510 262989
rect 298200 254175 298510 262961
rect 298200 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298510 254175
rect 298200 254113 298510 254147
rect 298200 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298510 254113
rect 298200 254051 298510 254085
rect 298200 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298510 254051
rect 298200 253989 298510 254023
rect 298200 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298510 253989
rect 298200 245175 298510 253961
rect 298200 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298510 245175
rect 298200 245113 298510 245147
rect 298200 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298510 245113
rect 298200 245051 298510 245085
rect 298200 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298510 245051
rect 298200 244989 298510 245023
rect 298200 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298510 244989
rect 298200 236175 298510 244961
rect 298200 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298510 236175
rect 298200 236113 298510 236147
rect 298200 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298510 236113
rect 298200 236051 298510 236085
rect 298200 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298510 236051
rect 298200 235989 298510 236023
rect 298200 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298510 235989
rect 298200 227175 298510 235961
rect 298200 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298510 227175
rect 298200 227113 298510 227147
rect 298200 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298510 227113
rect 298200 227051 298510 227085
rect 298200 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298510 227051
rect 298200 226989 298510 227023
rect 298200 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298510 226989
rect 298200 218175 298510 226961
rect 298200 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298510 218175
rect 298200 218113 298510 218147
rect 298200 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298510 218113
rect 298200 218051 298510 218085
rect 298200 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298510 218051
rect 298200 217989 298510 218023
rect 298200 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298510 217989
rect 298200 209175 298510 217961
rect 298200 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298510 209175
rect 298200 209113 298510 209147
rect 298200 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298510 209113
rect 298200 209051 298510 209085
rect 298200 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298510 209051
rect 298200 208989 298510 209023
rect 298200 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298510 208989
rect 298200 200175 298510 208961
rect 298200 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298510 200175
rect 298200 200113 298510 200147
rect 298200 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298510 200113
rect 298200 200051 298510 200085
rect 298200 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298510 200051
rect 298200 199989 298510 200023
rect 298200 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298510 199989
rect 298200 191175 298510 199961
rect 298200 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298510 191175
rect 298200 191113 298510 191147
rect 298200 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298510 191113
rect 298200 191051 298510 191085
rect 298200 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298510 191051
rect 298200 190989 298510 191023
rect 298200 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298510 190989
rect 298200 182175 298510 190961
rect 298200 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298510 182175
rect 298200 182113 298510 182147
rect 298200 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298510 182113
rect 298200 182051 298510 182085
rect 298200 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298510 182051
rect 298200 181989 298510 182023
rect 298200 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298510 181989
rect 298200 173175 298510 181961
rect 298200 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298510 173175
rect 298200 173113 298510 173147
rect 298200 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298510 173113
rect 298200 173051 298510 173085
rect 298200 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298510 173051
rect 298200 172989 298510 173023
rect 298200 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298510 172989
rect 298200 164175 298510 172961
rect 298200 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298510 164175
rect 298200 164113 298510 164147
rect 298200 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298510 164113
rect 298200 164051 298510 164085
rect 298200 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298510 164051
rect 298200 163989 298510 164023
rect 298200 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298510 163989
rect 298200 155175 298510 163961
rect 298200 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298510 155175
rect 298200 155113 298510 155147
rect 298200 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298510 155113
rect 298200 155051 298510 155085
rect 298200 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298510 155051
rect 298200 154989 298510 155023
rect 298200 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298510 154989
rect 298200 146175 298510 154961
rect 298200 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298510 146175
rect 298200 146113 298510 146147
rect 298200 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298510 146113
rect 298200 146051 298510 146085
rect 298200 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298510 146051
rect 298200 145989 298510 146023
rect 298200 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298510 145989
rect 298200 137175 298510 145961
rect 298200 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298510 137175
rect 298200 137113 298510 137147
rect 298200 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298510 137113
rect 298200 137051 298510 137085
rect 298200 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298510 137051
rect 298200 136989 298510 137023
rect 298200 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298510 136989
rect 298200 128175 298510 136961
rect 298200 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298510 128175
rect 298200 128113 298510 128147
rect 298200 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298510 128113
rect 298200 128051 298510 128085
rect 298200 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298510 128051
rect 298200 127989 298510 128023
rect 298200 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298510 127989
rect 298200 119175 298510 127961
rect 298200 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298510 119175
rect 298200 119113 298510 119147
rect 298200 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298510 119113
rect 298200 119051 298510 119085
rect 298200 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298510 119051
rect 298200 118989 298510 119023
rect 298200 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298510 118989
rect 298200 110175 298510 118961
rect 298200 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298510 110175
rect 298200 110113 298510 110147
rect 298200 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298510 110113
rect 298200 110051 298510 110085
rect 298200 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298510 110051
rect 298200 109989 298510 110023
rect 298200 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298510 109989
rect 298200 101175 298510 109961
rect 298200 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298510 101175
rect 298200 101113 298510 101147
rect 298200 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298510 101113
rect 298200 101051 298510 101085
rect 298200 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298510 101051
rect 298200 100989 298510 101023
rect 298200 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298510 100989
rect 298200 92175 298510 100961
rect 298200 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298510 92175
rect 298200 92113 298510 92147
rect 298200 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298510 92113
rect 298200 92051 298510 92085
rect 298200 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298510 92051
rect 298200 91989 298510 92023
rect 298200 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298510 91989
rect 298200 83175 298510 91961
rect 298200 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298510 83175
rect 298200 83113 298510 83147
rect 298200 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298510 83113
rect 298200 83051 298510 83085
rect 298200 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298510 83051
rect 298200 82989 298510 83023
rect 298200 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298510 82989
rect 298200 74175 298510 82961
rect 298200 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298510 74175
rect 298200 74113 298510 74147
rect 298200 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298510 74113
rect 298200 74051 298510 74085
rect 298200 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298510 74051
rect 298200 73989 298510 74023
rect 298200 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298510 73989
rect 298200 65175 298510 73961
rect 298200 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298510 65175
rect 298200 65113 298510 65147
rect 298200 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298510 65113
rect 298200 65051 298510 65085
rect 298200 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298510 65051
rect 298200 64989 298510 65023
rect 298200 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298510 64989
rect 298200 56175 298510 64961
rect 298200 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298510 56175
rect 298200 56113 298510 56147
rect 298200 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298510 56113
rect 298200 56051 298510 56085
rect 298200 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298510 56051
rect 298200 55989 298510 56023
rect 298200 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298510 55989
rect 298200 47175 298510 55961
rect 298200 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298510 47175
rect 298200 47113 298510 47147
rect 298200 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298510 47113
rect 298200 47051 298510 47085
rect 298200 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298510 47051
rect 298200 46989 298510 47023
rect 298200 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298510 46989
rect 298200 38175 298510 46961
rect 298200 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298510 38175
rect 298200 38113 298510 38147
rect 298200 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298510 38113
rect 298200 38051 298510 38085
rect 298200 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298510 38051
rect 298200 37989 298510 38023
rect 298200 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298510 37989
rect 298200 29175 298510 37961
rect 298200 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298510 29175
rect 298200 29113 298510 29147
rect 298200 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298510 29113
rect 298200 29051 298510 29085
rect 298200 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298510 29051
rect 298200 28989 298510 29023
rect 298200 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298510 28989
rect 298200 20175 298510 28961
rect 298200 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298510 20175
rect 298200 20113 298510 20147
rect 298200 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298510 20113
rect 298200 20051 298510 20085
rect 298200 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298510 20051
rect 298200 19989 298510 20023
rect 298200 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298510 19989
rect 298200 11175 298510 19961
rect 298200 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298510 11175
rect 298200 11113 298510 11147
rect 298200 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298510 11113
rect 298200 11051 298510 11085
rect 298200 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298510 11051
rect 298200 10989 298510 11023
rect 298200 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298510 10989
rect 298200 2175 298510 10961
rect 298200 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298510 2175
rect 298200 2113 298510 2147
rect 298200 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298510 2113
rect 298200 2051 298510 2085
rect 298200 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298510 2051
rect 298200 1989 298510 2023
rect 298200 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298510 1989
rect 298200 -80 298510 1961
rect 298200 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect 298200 -142 298510 -108
rect 298200 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect 298200 -204 298510 -170
rect 298200 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect 298200 -266 298510 -232
rect 298200 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect 298200 -342 298510 -294
rect 298680 293175 298990 298872
rect 298680 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect 298680 293113 298990 293147
rect 298680 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect 298680 293051 298990 293085
rect 298680 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect 298680 292989 298990 293023
rect 298680 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect 298680 284175 298990 292961
rect 298680 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect 298680 284113 298990 284147
rect 298680 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect 298680 284051 298990 284085
rect 298680 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect 298680 283989 298990 284023
rect 298680 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect 298680 275175 298990 283961
rect 298680 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect 298680 275113 298990 275147
rect 298680 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect 298680 275051 298990 275085
rect 298680 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect 298680 274989 298990 275023
rect 298680 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect 298680 266175 298990 274961
rect 298680 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect 298680 266113 298990 266147
rect 298680 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect 298680 266051 298990 266085
rect 298680 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect 298680 265989 298990 266023
rect 298680 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect 298680 257175 298990 265961
rect 298680 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect 298680 257113 298990 257147
rect 298680 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect 298680 257051 298990 257085
rect 298680 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect 298680 256989 298990 257023
rect 298680 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect 298680 248175 298990 256961
rect 298680 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect 298680 248113 298990 248147
rect 298680 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect 298680 248051 298990 248085
rect 298680 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect 298680 247989 298990 248023
rect 298680 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect 298680 239175 298990 247961
rect 298680 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect 298680 239113 298990 239147
rect 298680 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect 298680 239051 298990 239085
rect 298680 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect 298680 238989 298990 239023
rect 298680 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect 298680 230175 298990 238961
rect 298680 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect 298680 230113 298990 230147
rect 298680 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect 298680 230051 298990 230085
rect 298680 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect 298680 229989 298990 230023
rect 298680 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect 298680 221175 298990 229961
rect 298680 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect 298680 221113 298990 221147
rect 298680 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect 298680 221051 298990 221085
rect 298680 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect 298680 220989 298990 221023
rect 298680 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect 298680 212175 298990 220961
rect 298680 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect 298680 212113 298990 212147
rect 298680 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect 298680 212051 298990 212085
rect 298680 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect 298680 211989 298990 212023
rect 298680 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect 298680 203175 298990 211961
rect 298680 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect 298680 203113 298990 203147
rect 298680 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect 298680 203051 298990 203085
rect 298680 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect 298680 202989 298990 203023
rect 298680 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect 298680 194175 298990 202961
rect 298680 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect 298680 194113 298990 194147
rect 298680 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect 298680 194051 298990 194085
rect 298680 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect 298680 193989 298990 194023
rect 298680 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect 298680 185175 298990 193961
rect 298680 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect 298680 185113 298990 185147
rect 298680 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect 298680 185051 298990 185085
rect 298680 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect 298680 184989 298990 185023
rect 298680 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect 298680 176175 298990 184961
rect 298680 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect 298680 176113 298990 176147
rect 298680 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect 298680 176051 298990 176085
rect 298680 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect 298680 175989 298990 176023
rect 298680 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect 298680 167175 298990 175961
rect 298680 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect 298680 167113 298990 167147
rect 298680 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect 298680 167051 298990 167085
rect 298680 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect 298680 166989 298990 167023
rect 298680 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect 298680 158175 298990 166961
rect 298680 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect 298680 158113 298990 158147
rect 298680 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect 298680 158051 298990 158085
rect 298680 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect 298680 157989 298990 158023
rect 298680 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect 298680 149175 298990 157961
rect 298680 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect 298680 149113 298990 149147
rect 298680 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect 298680 149051 298990 149085
rect 298680 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect 298680 148989 298990 149023
rect 298680 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect 298680 140175 298990 148961
rect 298680 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect 298680 140113 298990 140147
rect 298680 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect 298680 140051 298990 140085
rect 298680 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect 298680 139989 298990 140023
rect 298680 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect 298680 131175 298990 139961
rect 298680 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect 298680 131113 298990 131147
rect 298680 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect 298680 131051 298990 131085
rect 298680 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect 298680 130989 298990 131023
rect 298680 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect 298680 122175 298990 130961
rect 298680 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect 298680 122113 298990 122147
rect 298680 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect 298680 122051 298990 122085
rect 298680 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect 298680 121989 298990 122023
rect 298680 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect 298680 113175 298990 121961
rect 298680 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect 298680 113113 298990 113147
rect 298680 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect 298680 113051 298990 113085
rect 298680 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect 298680 112989 298990 113023
rect 298680 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect 298680 104175 298990 112961
rect 298680 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect 298680 104113 298990 104147
rect 298680 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect 298680 104051 298990 104085
rect 298680 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect 298680 103989 298990 104023
rect 298680 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect 298680 95175 298990 103961
rect 298680 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect 298680 95113 298990 95147
rect 298680 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect 298680 95051 298990 95085
rect 298680 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect 298680 94989 298990 95023
rect 298680 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect 298680 86175 298990 94961
rect 298680 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect 298680 86113 298990 86147
rect 298680 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect 298680 86051 298990 86085
rect 298680 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect 298680 85989 298990 86023
rect 298680 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect 298680 77175 298990 85961
rect 298680 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect 298680 77113 298990 77147
rect 298680 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect 298680 77051 298990 77085
rect 298680 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect 298680 76989 298990 77023
rect 298680 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect 298680 68175 298990 76961
rect 298680 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect 298680 68113 298990 68147
rect 298680 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect 298680 68051 298990 68085
rect 298680 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect 298680 67989 298990 68023
rect 298680 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect 298680 59175 298990 67961
rect 298680 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect 298680 59113 298990 59147
rect 298680 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect 298680 59051 298990 59085
rect 298680 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect 298680 58989 298990 59023
rect 298680 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect 298680 50175 298990 58961
rect 298680 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect 298680 50113 298990 50147
rect 298680 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect 298680 50051 298990 50085
rect 298680 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect 298680 49989 298990 50023
rect 298680 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect 298680 41175 298990 49961
rect 298680 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect 298680 41113 298990 41147
rect 298680 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect 298680 41051 298990 41085
rect 298680 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect 298680 40989 298990 41023
rect 298680 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect 298680 32175 298990 40961
rect 298680 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect 298680 32113 298990 32147
rect 298680 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect 298680 32051 298990 32085
rect 298680 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect 298680 31989 298990 32023
rect 298680 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect 298680 23175 298990 31961
rect 298680 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect 298680 23113 298990 23147
rect 298680 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect 298680 23051 298990 23085
rect 298680 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect 298680 22989 298990 23023
rect 298680 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect 298680 14175 298990 22961
rect 298680 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect 298680 14113 298990 14147
rect 298680 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect 298680 14051 298990 14085
rect 298680 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect 298680 13989 298990 14023
rect 298680 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect 298680 5175 298990 13961
rect 298680 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect 298680 5113 298990 5147
rect 298680 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect 298680 5051 298990 5085
rect 298680 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect 298680 4989 298990 5023
rect 298680 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect 296409 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 296719 -560
rect 296409 -622 296719 -588
rect 296409 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 296719 -622
rect 296409 -684 296719 -650
rect 296409 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 296719 -684
rect 296409 -746 296719 -712
rect 296409 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 296719 -746
rect 296409 -822 296719 -774
rect 298680 -560 298990 4961
rect 298680 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect 298680 -622 298990 -588
rect 298680 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect 298680 -684 298990 -650
rect 298680 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect 298680 -746 298990 -712
rect 298680 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect 298680 -822 298990 -774
<< via4 >>
rect -910 299058 -882 299086
rect -848 299058 -820 299086
rect -786 299058 -758 299086
rect -724 299058 -696 299086
rect -910 298996 -882 299024
rect -848 298996 -820 299024
rect -786 298996 -758 299024
rect -724 298996 -696 299024
rect -910 298934 -882 298962
rect -848 298934 -820 298962
rect -786 298934 -758 298962
rect -724 298934 -696 298962
rect -910 298872 -882 298900
rect -848 298872 -820 298900
rect -786 298872 -758 298900
rect -724 298872 -696 298900
rect -910 293147 -882 293175
rect -848 293147 -820 293175
rect -786 293147 -758 293175
rect -724 293147 -696 293175
rect -910 293085 -882 293113
rect -848 293085 -820 293113
rect -786 293085 -758 293113
rect -724 293085 -696 293113
rect -910 293023 -882 293051
rect -848 293023 -820 293051
rect -786 293023 -758 293051
rect -724 293023 -696 293051
rect -910 292961 -882 292989
rect -848 292961 -820 292989
rect -786 292961 -758 292989
rect -724 292961 -696 292989
rect -910 284147 -882 284175
rect -848 284147 -820 284175
rect -786 284147 -758 284175
rect -724 284147 -696 284175
rect -910 284085 -882 284113
rect -848 284085 -820 284113
rect -786 284085 -758 284113
rect -724 284085 -696 284113
rect -910 284023 -882 284051
rect -848 284023 -820 284051
rect -786 284023 -758 284051
rect -724 284023 -696 284051
rect -910 283961 -882 283989
rect -848 283961 -820 283989
rect -786 283961 -758 283989
rect -724 283961 -696 283989
rect -910 275147 -882 275175
rect -848 275147 -820 275175
rect -786 275147 -758 275175
rect -724 275147 -696 275175
rect -910 275085 -882 275113
rect -848 275085 -820 275113
rect -786 275085 -758 275113
rect -724 275085 -696 275113
rect -910 275023 -882 275051
rect -848 275023 -820 275051
rect -786 275023 -758 275051
rect -724 275023 -696 275051
rect -910 274961 -882 274989
rect -848 274961 -820 274989
rect -786 274961 -758 274989
rect -724 274961 -696 274989
rect -910 266147 -882 266175
rect -848 266147 -820 266175
rect -786 266147 -758 266175
rect -724 266147 -696 266175
rect -910 266085 -882 266113
rect -848 266085 -820 266113
rect -786 266085 -758 266113
rect -724 266085 -696 266113
rect -910 266023 -882 266051
rect -848 266023 -820 266051
rect -786 266023 -758 266051
rect -724 266023 -696 266051
rect -910 265961 -882 265989
rect -848 265961 -820 265989
rect -786 265961 -758 265989
rect -724 265961 -696 265989
rect -910 257147 -882 257175
rect -848 257147 -820 257175
rect -786 257147 -758 257175
rect -724 257147 -696 257175
rect -910 257085 -882 257113
rect -848 257085 -820 257113
rect -786 257085 -758 257113
rect -724 257085 -696 257113
rect -910 257023 -882 257051
rect -848 257023 -820 257051
rect -786 257023 -758 257051
rect -724 257023 -696 257051
rect -910 256961 -882 256989
rect -848 256961 -820 256989
rect -786 256961 -758 256989
rect -724 256961 -696 256989
rect -910 248147 -882 248175
rect -848 248147 -820 248175
rect -786 248147 -758 248175
rect -724 248147 -696 248175
rect -910 248085 -882 248113
rect -848 248085 -820 248113
rect -786 248085 -758 248113
rect -724 248085 -696 248113
rect -910 248023 -882 248051
rect -848 248023 -820 248051
rect -786 248023 -758 248051
rect -724 248023 -696 248051
rect -910 247961 -882 247989
rect -848 247961 -820 247989
rect -786 247961 -758 247989
rect -724 247961 -696 247989
rect -910 239147 -882 239175
rect -848 239147 -820 239175
rect -786 239147 -758 239175
rect -724 239147 -696 239175
rect -910 239085 -882 239113
rect -848 239085 -820 239113
rect -786 239085 -758 239113
rect -724 239085 -696 239113
rect -910 239023 -882 239051
rect -848 239023 -820 239051
rect -786 239023 -758 239051
rect -724 239023 -696 239051
rect -910 238961 -882 238989
rect -848 238961 -820 238989
rect -786 238961 -758 238989
rect -724 238961 -696 238989
rect -910 230147 -882 230175
rect -848 230147 -820 230175
rect -786 230147 -758 230175
rect -724 230147 -696 230175
rect -910 230085 -882 230113
rect -848 230085 -820 230113
rect -786 230085 -758 230113
rect -724 230085 -696 230113
rect -910 230023 -882 230051
rect -848 230023 -820 230051
rect -786 230023 -758 230051
rect -724 230023 -696 230051
rect -910 229961 -882 229989
rect -848 229961 -820 229989
rect -786 229961 -758 229989
rect -724 229961 -696 229989
rect -910 221147 -882 221175
rect -848 221147 -820 221175
rect -786 221147 -758 221175
rect -724 221147 -696 221175
rect -910 221085 -882 221113
rect -848 221085 -820 221113
rect -786 221085 -758 221113
rect -724 221085 -696 221113
rect -910 221023 -882 221051
rect -848 221023 -820 221051
rect -786 221023 -758 221051
rect -724 221023 -696 221051
rect -910 220961 -882 220989
rect -848 220961 -820 220989
rect -786 220961 -758 220989
rect -724 220961 -696 220989
rect -910 212147 -882 212175
rect -848 212147 -820 212175
rect -786 212147 -758 212175
rect -724 212147 -696 212175
rect -910 212085 -882 212113
rect -848 212085 -820 212113
rect -786 212085 -758 212113
rect -724 212085 -696 212113
rect -910 212023 -882 212051
rect -848 212023 -820 212051
rect -786 212023 -758 212051
rect -724 212023 -696 212051
rect -910 211961 -882 211989
rect -848 211961 -820 211989
rect -786 211961 -758 211989
rect -724 211961 -696 211989
rect -910 203147 -882 203175
rect -848 203147 -820 203175
rect -786 203147 -758 203175
rect -724 203147 -696 203175
rect -910 203085 -882 203113
rect -848 203085 -820 203113
rect -786 203085 -758 203113
rect -724 203085 -696 203113
rect -910 203023 -882 203051
rect -848 203023 -820 203051
rect -786 203023 -758 203051
rect -724 203023 -696 203051
rect -910 202961 -882 202989
rect -848 202961 -820 202989
rect -786 202961 -758 202989
rect -724 202961 -696 202989
rect -910 194147 -882 194175
rect -848 194147 -820 194175
rect -786 194147 -758 194175
rect -724 194147 -696 194175
rect -910 194085 -882 194113
rect -848 194085 -820 194113
rect -786 194085 -758 194113
rect -724 194085 -696 194113
rect -910 194023 -882 194051
rect -848 194023 -820 194051
rect -786 194023 -758 194051
rect -724 194023 -696 194051
rect -910 193961 -882 193989
rect -848 193961 -820 193989
rect -786 193961 -758 193989
rect -724 193961 -696 193989
rect -910 185147 -882 185175
rect -848 185147 -820 185175
rect -786 185147 -758 185175
rect -724 185147 -696 185175
rect -910 185085 -882 185113
rect -848 185085 -820 185113
rect -786 185085 -758 185113
rect -724 185085 -696 185113
rect -910 185023 -882 185051
rect -848 185023 -820 185051
rect -786 185023 -758 185051
rect -724 185023 -696 185051
rect -910 184961 -882 184989
rect -848 184961 -820 184989
rect -786 184961 -758 184989
rect -724 184961 -696 184989
rect -910 176147 -882 176175
rect -848 176147 -820 176175
rect -786 176147 -758 176175
rect -724 176147 -696 176175
rect -910 176085 -882 176113
rect -848 176085 -820 176113
rect -786 176085 -758 176113
rect -724 176085 -696 176113
rect -910 176023 -882 176051
rect -848 176023 -820 176051
rect -786 176023 -758 176051
rect -724 176023 -696 176051
rect -910 175961 -882 175989
rect -848 175961 -820 175989
rect -786 175961 -758 175989
rect -724 175961 -696 175989
rect -910 167147 -882 167175
rect -848 167147 -820 167175
rect -786 167147 -758 167175
rect -724 167147 -696 167175
rect -910 167085 -882 167113
rect -848 167085 -820 167113
rect -786 167085 -758 167113
rect -724 167085 -696 167113
rect -910 167023 -882 167051
rect -848 167023 -820 167051
rect -786 167023 -758 167051
rect -724 167023 -696 167051
rect -910 166961 -882 166989
rect -848 166961 -820 166989
rect -786 166961 -758 166989
rect -724 166961 -696 166989
rect -910 158147 -882 158175
rect -848 158147 -820 158175
rect -786 158147 -758 158175
rect -724 158147 -696 158175
rect -910 158085 -882 158113
rect -848 158085 -820 158113
rect -786 158085 -758 158113
rect -724 158085 -696 158113
rect -910 158023 -882 158051
rect -848 158023 -820 158051
rect -786 158023 -758 158051
rect -724 158023 -696 158051
rect -910 157961 -882 157989
rect -848 157961 -820 157989
rect -786 157961 -758 157989
rect -724 157961 -696 157989
rect -910 149147 -882 149175
rect -848 149147 -820 149175
rect -786 149147 -758 149175
rect -724 149147 -696 149175
rect -910 149085 -882 149113
rect -848 149085 -820 149113
rect -786 149085 -758 149113
rect -724 149085 -696 149113
rect -910 149023 -882 149051
rect -848 149023 -820 149051
rect -786 149023 -758 149051
rect -724 149023 -696 149051
rect -910 148961 -882 148989
rect -848 148961 -820 148989
rect -786 148961 -758 148989
rect -724 148961 -696 148989
rect -910 140147 -882 140175
rect -848 140147 -820 140175
rect -786 140147 -758 140175
rect -724 140147 -696 140175
rect -910 140085 -882 140113
rect -848 140085 -820 140113
rect -786 140085 -758 140113
rect -724 140085 -696 140113
rect -910 140023 -882 140051
rect -848 140023 -820 140051
rect -786 140023 -758 140051
rect -724 140023 -696 140051
rect -910 139961 -882 139989
rect -848 139961 -820 139989
rect -786 139961 -758 139989
rect -724 139961 -696 139989
rect -910 131147 -882 131175
rect -848 131147 -820 131175
rect -786 131147 -758 131175
rect -724 131147 -696 131175
rect -910 131085 -882 131113
rect -848 131085 -820 131113
rect -786 131085 -758 131113
rect -724 131085 -696 131113
rect -910 131023 -882 131051
rect -848 131023 -820 131051
rect -786 131023 -758 131051
rect -724 131023 -696 131051
rect -910 130961 -882 130989
rect -848 130961 -820 130989
rect -786 130961 -758 130989
rect -724 130961 -696 130989
rect -910 122147 -882 122175
rect -848 122147 -820 122175
rect -786 122147 -758 122175
rect -724 122147 -696 122175
rect -910 122085 -882 122113
rect -848 122085 -820 122113
rect -786 122085 -758 122113
rect -724 122085 -696 122113
rect -910 122023 -882 122051
rect -848 122023 -820 122051
rect -786 122023 -758 122051
rect -724 122023 -696 122051
rect -910 121961 -882 121989
rect -848 121961 -820 121989
rect -786 121961 -758 121989
rect -724 121961 -696 121989
rect -910 113147 -882 113175
rect -848 113147 -820 113175
rect -786 113147 -758 113175
rect -724 113147 -696 113175
rect -910 113085 -882 113113
rect -848 113085 -820 113113
rect -786 113085 -758 113113
rect -724 113085 -696 113113
rect -910 113023 -882 113051
rect -848 113023 -820 113051
rect -786 113023 -758 113051
rect -724 113023 -696 113051
rect -910 112961 -882 112989
rect -848 112961 -820 112989
rect -786 112961 -758 112989
rect -724 112961 -696 112989
rect -910 104147 -882 104175
rect -848 104147 -820 104175
rect -786 104147 -758 104175
rect -724 104147 -696 104175
rect -910 104085 -882 104113
rect -848 104085 -820 104113
rect -786 104085 -758 104113
rect -724 104085 -696 104113
rect -910 104023 -882 104051
rect -848 104023 -820 104051
rect -786 104023 -758 104051
rect -724 104023 -696 104051
rect -910 103961 -882 103989
rect -848 103961 -820 103989
rect -786 103961 -758 103989
rect -724 103961 -696 103989
rect -910 95147 -882 95175
rect -848 95147 -820 95175
rect -786 95147 -758 95175
rect -724 95147 -696 95175
rect -910 95085 -882 95113
rect -848 95085 -820 95113
rect -786 95085 -758 95113
rect -724 95085 -696 95113
rect -910 95023 -882 95051
rect -848 95023 -820 95051
rect -786 95023 -758 95051
rect -724 95023 -696 95051
rect -910 94961 -882 94989
rect -848 94961 -820 94989
rect -786 94961 -758 94989
rect -724 94961 -696 94989
rect -910 86147 -882 86175
rect -848 86147 -820 86175
rect -786 86147 -758 86175
rect -724 86147 -696 86175
rect -910 86085 -882 86113
rect -848 86085 -820 86113
rect -786 86085 -758 86113
rect -724 86085 -696 86113
rect -910 86023 -882 86051
rect -848 86023 -820 86051
rect -786 86023 -758 86051
rect -724 86023 -696 86051
rect -910 85961 -882 85989
rect -848 85961 -820 85989
rect -786 85961 -758 85989
rect -724 85961 -696 85989
rect -910 77147 -882 77175
rect -848 77147 -820 77175
rect -786 77147 -758 77175
rect -724 77147 -696 77175
rect -910 77085 -882 77113
rect -848 77085 -820 77113
rect -786 77085 -758 77113
rect -724 77085 -696 77113
rect -910 77023 -882 77051
rect -848 77023 -820 77051
rect -786 77023 -758 77051
rect -724 77023 -696 77051
rect -910 76961 -882 76989
rect -848 76961 -820 76989
rect -786 76961 -758 76989
rect -724 76961 -696 76989
rect -910 68147 -882 68175
rect -848 68147 -820 68175
rect -786 68147 -758 68175
rect -724 68147 -696 68175
rect -910 68085 -882 68113
rect -848 68085 -820 68113
rect -786 68085 -758 68113
rect -724 68085 -696 68113
rect -910 68023 -882 68051
rect -848 68023 -820 68051
rect -786 68023 -758 68051
rect -724 68023 -696 68051
rect -910 67961 -882 67989
rect -848 67961 -820 67989
rect -786 67961 -758 67989
rect -724 67961 -696 67989
rect -910 59147 -882 59175
rect -848 59147 -820 59175
rect -786 59147 -758 59175
rect -724 59147 -696 59175
rect -910 59085 -882 59113
rect -848 59085 -820 59113
rect -786 59085 -758 59113
rect -724 59085 -696 59113
rect -910 59023 -882 59051
rect -848 59023 -820 59051
rect -786 59023 -758 59051
rect -724 59023 -696 59051
rect -910 58961 -882 58989
rect -848 58961 -820 58989
rect -786 58961 -758 58989
rect -724 58961 -696 58989
rect -910 50147 -882 50175
rect -848 50147 -820 50175
rect -786 50147 -758 50175
rect -724 50147 -696 50175
rect -910 50085 -882 50113
rect -848 50085 -820 50113
rect -786 50085 -758 50113
rect -724 50085 -696 50113
rect -910 50023 -882 50051
rect -848 50023 -820 50051
rect -786 50023 -758 50051
rect -724 50023 -696 50051
rect -910 49961 -882 49989
rect -848 49961 -820 49989
rect -786 49961 -758 49989
rect -724 49961 -696 49989
rect -910 41147 -882 41175
rect -848 41147 -820 41175
rect -786 41147 -758 41175
rect -724 41147 -696 41175
rect -910 41085 -882 41113
rect -848 41085 -820 41113
rect -786 41085 -758 41113
rect -724 41085 -696 41113
rect -910 41023 -882 41051
rect -848 41023 -820 41051
rect -786 41023 -758 41051
rect -724 41023 -696 41051
rect -910 40961 -882 40989
rect -848 40961 -820 40989
rect -786 40961 -758 40989
rect -724 40961 -696 40989
rect -910 32147 -882 32175
rect -848 32147 -820 32175
rect -786 32147 -758 32175
rect -724 32147 -696 32175
rect -910 32085 -882 32113
rect -848 32085 -820 32113
rect -786 32085 -758 32113
rect -724 32085 -696 32113
rect -910 32023 -882 32051
rect -848 32023 -820 32051
rect -786 32023 -758 32051
rect -724 32023 -696 32051
rect -910 31961 -882 31989
rect -848 31961 -820 31989
rect -786 31961 -758 31989
rect -724 31961 -696 31989
rect -910 23147 -882 23175
rect -848 23147 -820 23175
rect -786 23147 -758 23175
rect -724 23147 -696 23175
rect -910 23085 -882 23113
rect -848 23085 -820 23113
rect -786 23085 -758 23113
rect -724 23085 -696 23113
rect -910 23023 -882 23051
rect -848 23023 -820 23051
rect -786 23023 -758 23051
rect -724 23023 -696 23051
rect -910 22961 -882 22989
rect -848 22961 -820 22989
rect -786 22961 -758 22989
rect -724 22961 -696 22989
rect -910 14147 -882 14175
rect -848 14147 -820 14175
rect -786 14147 -758 14175
rect -724 14147 -696 14175
rect -910 14085 -882 14113
rect -848 14085 -820 14113
rect -786 14085 -758 14113
rect -724 14085 -696 14113
rect -910 14023 -882 14051
rect -848 14023 -820 14051
rect -786 14023 -758 14051
rect -724 14023 -696 14051
rect -910 13961 -882 13989
rect -848 13961 -820 13989
rect -786 13961 -758 13989
rect -724 13961 -696 13989
rect -910 5147 -882 5175
rect -848 5147 -820 5175
rect -786 5147 -758 5175
rect -724 5147 -696 5175
rect -910 5085 -882 5113
rect -848 5085 -820 5113
rect -786 5085 -758 5113
rect -724 5085 -696 5113
rect -910 5023 -882 5051
rect -848 5023 -820 5051
rect -786 5023 -758 5051
rect -724 5023 -696 5051
rect -910 4961 -882 4989
rect -848 4961 -820 4989
rect -786 4961 -758 4989
rect -724 4961 -696 4989
rect -430 298578 -402 298606
rect -368 298578 -340 298606
rect -306 298578 -278 298606
rect -244 298578 -216 298606
rect -430 298516 -402 298544
rect -368 298516 -340 298544
rect -306 298516 -278 298544
rect -244 298516 -216 298544
rect -430 298454 -402 298482
rect -368 298454 -340 298482
rect -306 298454 -278 298482
rect -244 298454 -216 298482
rect -430 298392 -402 298420
rect -368 298392 -340 298420
rect -306 298392 -278 298420
rect -244 298392 -216 298420
rect -430 290147 -402 290175
rect -368 290147 -340 290175
rect -306 290147 -278 290175
rect -244 290147 -216 290175
rect -430 290085 -402 290113
rect -368 290085 -340 290113
rect -306 290085 -278 290113
rect -244 290085 -216 290113
rect -430 290023 -402 290051
rect -368 290023 -340 290051
rect -306 290023 -278 290051
rect -244 290023 -216 290051
rect -430 289961 -402 289989
rect -368 289961 -340 289989
rect -306 289961 -278 289989
rect -244 289961 -216 289989
rect -430 281147 -402 281175
rect -368 281147 -340 281175
rect -306 281147 -278 281175
rect -244 281147 -216 281175
rect -430 281085 -402 281113
rect -368 281085 -340 281113
rect -306 281085 -278 281113
rect -244 281085 -216 281113
rect -430 281023 -402 281051
rect -368 281023 -340 281051
rect -306 281023 -278 281051
rect -244 281023 -216 281051
rect -430 280961 -402 280989
rect -368 280961 -340 280989
rect -306 280961 -278 280989
rect -244 280961 -216 280989
rect -430 272147 -402 272175
rect -368 272147 -340 272175
rect -306 272147 -278 272175
rect -244 272147 -216 272175
rect -430 272085 -402 272113
rect -368 272085 -340 272113
rect -306 272085 -278 272113
rect -244 272085 -216 272113
rect -430 272023 -402 272051
rect -368 272023 -340 272051
rect -306 272023 -278 272051
rect -244 272023 -216 272051
rect -430 271961 -402 271989
rect -368 271961 -340 271989
rect -306 271961 -278 271989
rect -244 271961 -216 271989
rect 2757 298578 2785 298606
rect 2819 298578 2847 298606
rect 2881 298578 2909 298606
rect 2943 298578 2971 298606
rect 2757 298516 2785 298544
rect 2819 298516 2847 298544
rect 2881 298516 2909 298544
rect 2943 298516 2971 298544
rect 2757 298454 2785 298482
rect 2819 298454 2847 298482
rect 2881 298454 2909 298482
rect 2943 298454 2971 298482
rect 2757 298392 2785 298420
rect 2819 298392 2847 298420
rect 2881 298392 2909 298420
rect 2943 298392 2971 298420
rect 2757 290147 2785 290175
rect 2819 290147 2847 290175
rect 2881 290147 2909 290175
rect 2943 290147 2971 290175
rect 2757 290085 2785 290113
rect 2819 290085 2847 290113
rect 2881 290085 2909 290113
rect 2943 290085 2971 290113
rect 2757 290023 2785 290051
rect 2819 290023 2847 290051
rect 2881 290023 2909 290051
rect 2943 290023 2971 290051
rect 2757 289961 2785 289989
rect 2819 289961 2847 289989
rect 2881 289961 2909 289989
rect 2943 289961 2971 289989
rect 2757 281147 2785 281175
rect 2819 281147 2847 281175
rect 2881 281147 2909 281175
rect 2943 281147 2971 281175
rect 2757 281085 2785 281113
rect 2819 281085 2847 281113
rect 2881 281085 2909 281113
rect 2943 281085 2971 281113
rect 2757 281023 2785 281051
rect 2819 281023 2847 281051
rect 2881 281023 2909 281051
rect 2943 281023 2971 281051
rect 2757 280961 2785 280989
rect 2819 280961 2847 280989
rect 2881 280961 2909 280989
rect 2943 280961 2971 280989
rect 2757 272147 2785 272175
rect 2819 272147 2847 272175
rect 2881 272147 2909 272175
rect 2943 272147 2971 272175
rect 2757 272085 2785 272113
rect 2819 272085 2847 272113
rect 2881 272085 2909 272113
rect 2943 272085 2971 272113
rect 2757 272023 2785 272051
rect 2819 272023 2847 272051
rect 2881 272023 2909 272051
rect 2943 272023 2971 272051
rect 2757 271961 2785 271989
rect 2819 271961 2847 271989
rect 2881 271961 2909 271989
rect 2943 271961 2971 271989
rect -430 263147 -402 263175
rect -368 263147 -340 263175
rect -306 263147 -278 263175
rect -244 263147 -216 263175
rect -430 263085 -402 263113
rect -368 263085 -340 263113
rect -306 263085 -278 263113
rect -244 263085 -216 263113
rect -430 263023 -402 263051
rect -368 263023 -340 263051
rect -306 263023 -278 263051
rect -244 263023 -216 263051
rect -430 262961 -402 262989
rect -368 262961 -340 262989
rect -306 262961 -278 262989
rect -244 262961 -216 262989
rect -430 254147 -402 254175
rect -368 254147 -340 254175
rect -306 254147 -278 254175
rect -244 254147 -216 254175
rect -430 254085 -402 254113
rect -368 254085 -340 254113
rect -306 254085 -278 254113
rect -244 254085 -216 254113
rect -430 254023 -402 254051
rect -368 254023 -340 254051
rect -306 254023 -278 254051
rect -244 254023 -216 254051
rect -430 253961 -402 253989
rect -368 253961 -340 253989
rect -306 253961 -278 253989
rect -244 253961 -216 253989
rect -430 245147 -402 245175
rect -368 245147 -340 245175
rect -306 245147 -278 245175
rect -244 245147 -216 245175
rect -430 245085 -402 245113
rect -368 245085 -340 245113
rect -306 245085 -278 245113
rect -244 245085 -216 245113
rect -430 245023 -402 245051
rect -368 245023 -340 245051
rect -306 245023 -278 245051
rect -244 245023 -216 245051
rect -430 244961 -402 244989
rect -368 244961 -340 244989
rect -306 244961 -278 244989
rect -244 244961 -216 244989
rect -430 236147 -402 236175
rect -368 236147 -340 236175
rect -306 236147 -278 236175
rect -244 236147 -216 236175
rect -430 236085 -402 236113
rect -368 236085 -340 236113
rect -306 236085 -278 236113
rect -244 236085 -216 236113
rect -430 236023 -402 236051
rect -368 236023 -340 236051
rect -306 236023 -278 236051
rect -244 236023 -216 236051
rect -430 235961 -402 235989
rect -368 235961 -340 235989
rect -306 235961 -278 235989
rect -244 235961 -216 235989
rect -430 227147 -402 227175
rect -368 227147 -340 227175
rect -306 227147 -278 227175
rect -244 227147 -216 227175
rect -430 227085 -402 227113
rect -368 227085 -340 227113
rect -306 227085 -278 227113
rect -244 227085 -216 227113
rect -430 227023 -402 227051
rect -368 227023 -340 227051
rect -306 227023 -278 227051
rect -244 227023 -216 227051
rect -430 226961 -402 226989
rect -368 226961 -340 226989
rect -306 226961 -278 226989
rect -244 226961 -216 226989
rect -430 218147 -402 218175
rect -368 218147 -340 218175
rect -306 218147 -278 218175
rect -244 218147 -216 218175
rect -430 218085 -402 218113
rect -368 218085 -340 218113
rect -306 218085 -278 218113
rect -244 218085 -216 218113
rect -430 218023 -402 218051
rect -368 218023 -340 218051
rect -306 218023 -278 218051
rect -244 218023 -216 218051
rect -430 217961 -402 217989
rect -368 217961 -340 217989
rect -306 217961 -278 217989
rect -244 217961 -216 217989
rect -430 209147 -402 209175
rect -368 209147 -340 209175
rect -306 209147 -278 209175
rect -244 209147 -216 209175
rect -430 209085 -402 209113
rect -368 209085 -340 209113
rect -306 209085 -278 209113
rect -244 209085 -216 209113
rect -430 209023 -402 209051
rect -368 209023 -340 209051
rect -306 209023 -278 209051
rect -244 209023 -216 209051
rect -430 208961 -402 208989
rect -368 208961 -340 208989
rect -306 208961 -278 208989
rect -244 208961 -216 208989
rect -430 200147 -402 200175
rect -368 200147 -340 200175
rect -306 200147 -278 200175
rect -244 200147 -216 200175
rect -430 200085 -402 200113
rect -368 200085 -340 200113
rect -306 200085 -278 200113
rect -244 200085 -216 200113
rect -430 200023 -402 200051
rect -368 200023 -340 200051
rect -306 200023 -278 200051
rect -244 200023 -216 200051
rect -430 199961 -402 199989
rect -368 199961 -340 199989
rect -306 199961 -278 199989
rect -244 199961 -216 199989
rect -430 191147 -402 191175
rect -368 191147 -340 191175
rect -306 191147 -278 191175
rect -244 191147 -216 191175
rect -430 191085 -402 191113
rect -368 191085 -340 191113
rect -306 191085 -278 191113
rect -244 191085 -216 191113
rect -430 191023 -402 191051
rect -368 191023 -340 191051
rect -306 191023 -278 191051
rect -244 191023 -216 191051
rect -430 190961 -402 190989
rect -368 190961 -340 190989
rect -306 190961 -278 190989
rect -244 190961 -216 190989
rect -430 182147 -402 182175
rect -368 182147 -340 182175
rect -306 182147 -278 182175
rect -244 182147 -216 182175
rect -430 182085 -402 182113
rect -368 182085 -340 182113
rect -306 182085 -278 182113
rect -244 182085 -216 182113
rect -430 182023 -402 182051
rect -368 182023 -340 182051
rect -306 182023 -278 182051
rect -244 182023 -216 182051
rect -430 181961 -402 181989
rect -368 181961 -340 181989
rect -306 181961 -278 181989
rect -244 181961 -216 181989
rect -430 173147 -402 173175
rect -368 173147 -340 173175
rect -306 173147 -278 173175
rect -244 173147 -216 173175
rect -430 173085 -402 173113
rect -368 173085 -340 173113
rect -306 173085 -278 173113
rect -244 173085 -216 173113
rect -430 173023 -402 173051
rect -368 173023 -340 173051
rect -306 173023 -278 173051
rect -244 173023 -216 173051
rect -430 172961 -402 172989
rect -368 172961 -340 172989
rect -306 172961 -278 172989
rect -244 172961 -216 172989
rect -430 164147 -402 164175
rect -368 164147 -340 164175
rect -306 164147 -278 164175
rect -244 164147 -216 164175
rect -430 164085 -402 164113
rect -368 164085 -340 164113
rect -306 164085 -278 164113
rect -244 164085 -216 164113
rect -430 164023 -402 164051
rect -368 164023 -340 164051
rect -306 164023 -278 164051
rect -244 164023 -216 164051
rect -430 163961 -402 163989
rect -368 163961 -340 163989
rect -306 163961 -278 163989
rect -244 163961 -216 163989
rect 2757 263147 2785 263175
rect 2819 263147 2847 263175
rect 2881 263147 2909 263175
rect 2943 263147 2971 263175
rect 2757 263085 2785 263113
rect 2819 263085 2847 263113
rect 2881 263085 2909 263113
rect 2943 263085 2971 263113
rect 2757 263023 2785 263051
rect 2819 263023 2847 263051
rect 2881 263023 2909 263051
rect 2943 263023 2971 263051
rect 2757 262961 2785 262989
rect 2819 262961 2847 262989
rect 2881 262961 2909 262989
rect 2943 262961 2971 262989
rect 2757 254147 2785 254175
rect 2819 254147 2847 254175
rect 2881 254147 2909 254175
rect 2943 254147 2971 254175
rect 2757 254085 2785 254113
rect 2819 254085 2847 254113
rect 2881 254085 2909 254113
rect 2943 254085 2971 254113
rect 2757 254023 2785 254051
rect 2819 254023 2847 254051
rect 2881 254023 2909 254051
rect 2943 254023 2971 254051
rect 2757 253961 2785 253989
rect 2819 253961 2847 253989
rect 2881 253961 2909 253989
rect 2943 253961 2971 253989
rect -430 155147 -402 155175
rect -368 155147 -340 155175
rect -306 155147 -278 155175
rect -244 155147 -216 155175
rect -430 155085 -402 155113
rect -368 155085 -340 155113
rect -306 155085 -278 155113
rect -244 155085 -216 155113
rect -430 155023 -402 155051
rect -368 155023 -340 155051
rect -306 155023 -278 155051
rect -244 155023 -216 155051
rect -430 154961 -402 154989
rect -368 154961 -340 154989
rect -306 154961 -278 154989
rect -244 154961 -216 154989
rect -430 146147 -402 146175
rect -368 146147 -340 146175
rect -306 146147 -278 146175
rect -244 146147 -216 146175
rect -430 146085 -402 146113
rect -368 146085 -340 146113
rect -306 146085 -278 146113
rect -244 146085 -216 146113
rect -430 146023 -402 146051
rect -368 146023 -340 146051
rect -306 146023 -278 146051
rect -244 146023 -216 146051
rect -430 145961 -402 145989
rect -368 145961 -340 145989
rect -306 145961 -278 145989
rect -244 145961 -216 145989
rect -430 137147 -402 137175
rect -368 137147 -340 137175
rect -306 137147 -278 137175
rect -244 137147 -216 137175
rect -430 137085 -402 137113
rect -368 137085 -340 137113
rect -306 137085 -278 137113
rect -244 137085 -216 137113
rect -430 137023 -402 137051
rect -368 137023 -340 137051
rect -306 137023 -278 137051
rect -244 137023 -216 137051
rect -430 136961 -402 136989
rect -368 136961 -340 136989
rect -306 136961 -278 136989
rect -244 136961 -216 136989
rect -430 128147 -402 128175
rect -368 128147 -340 128175
rect -306 128147 -278 128175
rect -244 128147 -216 128175
rect -430 128085 -402 128113
rect -368 128085 -340 128113
rect -306 128085 -278 128113
rect -244 128085 -216 128113
rect -430 128023 -402 128051
rect -368 128023 -340 128051
rect -306 128023 -278 128051
rect -244 128023 -216 128051
rect -430 127961 -402 127989
rect -368 127961 -340 127989
rect -306 127961 -278 127989
rect -244 127961 -216 127989
rect -430 119147 -402 119175
rect -368 119147 -340 119175
rect -306 119147 -278 119175
rect -244 119147 -216 119175
rect -430 119085 -402 119113
rect -368 119085 -340 119113
rect -306 119085 -278 119113
rect -244 119085 -216 119113
rect -430 119023 -402 119051
rect -368 119023 -340 119051
rect -306 119023 -278 119051
rect -244 119023 -216 119051
rect -430 118961 -402 118989
rect -368 118961 -340 118989
rect -306 118961 -278 118989
rect -244 118961 -216 118989
rect -430 110147 -402 110175
rect -368 110147 -340 110175
rect -306 110147 -278 110175
rect -244 110147 -216 110175
rect -430 110085 -402 110113
rect -368 110085 -340 110113
rect -306 110085 -278 110113
rect -244 110085 -216 110113
rect -430 110023 -402 110051
rect -368 110023 -340 110051
rect -306 110023 -278 110051
rect -244 110023 -216 110051
rect -430 109961 -402 109989
rect -368 109961 -340 109989
rect -306 109961 -278 109989
rect -244 109961 -216 109989
rect -430 101147 -402 101175
rect -368 101147 -340 101175
rect -306 101147 -278 101175
rect -244 101147 -216 101175
rect -430 101085 -402 101113
rect -368 101085 -340 101113
rect -306 101085 -278 101113
rect -244 101085 -216 101113
rect -430 101023 -402 101051
rect -368 101023 -340 101051
rect -306 101023 -278 101051
rect -244 101023 -216 101051
rect -430 100961 -402 100989
rect -368 100961 -340 100989
rect -306 100961 -278 100989
rect -244 100961 -216 100989
rect -430 92147 -402 92175
rect -368 92147 -340 92175
rect -306 92147 -278 92175
rect -244 92147 -216 92175
rect -430 92085 -402 92113
rect -368 92085 -340 92113
rect -306 92085 -278 92113
rect -244 92085 -216 92113
rect -430 92023 -402 92051
rect -368 92023 -340 92051
rect -306 92023 -278 92051
rect -244 92023 -216 92051
rect -430 91961 -402 91989
rect -368 91961 -340 91989
rect -306 91961 -278 91989
rect -244 91961 -216 91989
rect -430 83147 -402 83175
rect -368 83147 -340 83175
rect -306 83147 -278 83175
rect -244 83147 -216 83175
rect -430 83085 -402 83113
rect -368 83085 -340 83113
rect -306 83085 -278 83113
rect -244 83085 -216 83113
rect -430 83023 -402 83051
rect -368 83023 -340 83051
rect -306 83023 -278 83051
rect -244 83023 -216 83051
rect -430 82961 -402 82989
rect -368 82961 -340 82989
rect -306 82961 -278 82989
rect -244 82961 -216 82989
rect -430 74147 -402 74175
rect -368 74147 -340 74175
rect -306 74147 -278 74175
rect -244 74147 -216 74175
rect -430 74085 -402 74113
rect -368 74085 -340 74113
rect -306 74085 -278 74113
rect -244 74085 -216 74113
rect -430 74023 -402 74051
rect -368 74023 -340 74051
rect -306 74023 -278 74051
rect -244 74023 -216 74051
rect -430 73961 -402 73989
rect -368 73961 -340 73989
rect -306 73961 -278 73989
rect -244 73961 -216 73989
rect -430 65147 -402 65175
rect -368 65147 -340 65175
rect -306 65147 -278 65175
rect -244 65147 -216 65175
rect -430 65085 -402 65113
rect -368 65085 -340 65113
rect -306 65085 -278 65113
rect -244 65085 -216 65113
rect -430 65023 -402 65051
rect -368 65023 -340 65051
rect -306 65023 -278 65051
rect -244 65023 -216 65051
rect -430 64961 -402 64989
rect -368 64961 -340 64989
rect -306 64961 -278 64989
rect -244 64961 -216 64989
rect -430 56147 -402 56175
rect -368 56147 -340 56175
rect -306 56147 -278 56175
rect -244 56147 -216 56175
rect -430 56085 -402 56113
rect -368 56085 -340 56113
rect -306 56085 -278 56113
rect -244 56085 -216 56113
rect -430 56023 -402 56051
rect -368 56023 -340 56051
rect -306 56023 -278 56051
rect -244 56023 -216 56051
rect -430 55961 -402 55989
rect -368 55961 -340 55989
rect -306 55961 -278 55989
rect -244 55961 -216 55989
rect 2757 245147 2785 245175
rect 2819 245147 2847 245175
rect 2881 245147 2909 245175
rect 2943 245147 2971 245175
rect 2757 245085 2785 245113
rect 2819 245085 2847 245113
rect 2881 245085 2909 245113
rect 2943 245085 2971 245113
rect 2757 245023 2785 245051
rect 2819 245023 2847 245051
rect 2881 245023 2909 245051
rect 2943 245023 2971 245051
rect 2757 244961 2785 244989
rect 2819 244961 2847 244989
rect 2881 244961 2909 244989
rect 2943 244961 2971 244989
rect 2757 236147 2785 236175
rect 2819 236147 2847 236175
rect 2881 236147 2909 236175
rect 2943 236147 2971 236175
rect 2757 236085 2785 236113
rect 2819 236085 2847 236113
rect 2881 236085 2909 236113
rect 2943 236085 2971 236113
rect 2757 236023 2785 236051
rect 2819 236023 2847 236051
rect 2881 236023 2909 236051
rect 2943 236023 2971 236051
rect 2757 235961 2785 235989
rect 2819 235961 2847 235989
rect 2881 235961 2909 235989
rect 2943 235961 2971 235989
rect 2757 227147 2785 227175
rect 2819 227147 2847 227175
rect 2881 227147 2909 227175
rect 2943 227147 2971 227175
rect 2757 227085 2785 227113
rect 2819 227085 2847 227113
rect 2881 227085 2909 227113
rect 2943 227085 2971 227113
rect 2757 227023 2785 227051
rect 2819 227023 2847 227051
rect 2881 227023 2909 227051
rect 2943 227023 2971 227051
rect 2757 226961 2785 226989
rect 2819 226961 2847 226989
rect 2881 226961 2909 226989
rect 2943 226961 2971 226989
rect -430 47147 -402 47175
rect -368 47147 -340 47175
rect -306 47147 -278 47175
rect -244 47147 -216 47175
rect -430 47085 -402 47113
rect -368 47085 -340 47113
rect -306 47085 -278 47113
rect -244 47085 -216 47113
rect -430 47023 -402 47051
rect -368 47023 -340 47051
rect -306 47023 -278 47051
rect -244 47023 -216 47051
rect -430 46961 -402 46989
rect -368 46961 -340 46989
rect -306 46961 -278 46989
rect -244 46961 -216 46989
rect -430 38147 -402 38175
rect -368 38147 -340 38175
rect -306 38147 -278 38175
rect -244 38147 -216 38175
rect -430 38085 -402 38113
rect -368 38085 -340 38113
rect -306 38085 -278 38113
rect -244 38085 -216 38113
rect -430 38023 -402 38051
rect -368 38023 -340 38051
rect -306 38023 -278 38051
rect -244 38023 -216 38051
rect -430 37961 -402 37989
rect -368 37961 -340 37989
rect -306 37961 -278 37989
rect -244 37961 -216 37989
rect 2757 218147 2785 218175
rect 2819 218147 2847 218175
rect 2881 218147 2909 218175
rect 2943 218147 2971 218175
rect 2757 218085 2785 218113
rect 2819 218085 2847 218113
rect 2881 218085 2909 218113
rect 2943 218085 2971 218113
rect 2757 218023 2785 218051
rect 2819 218023 2847 218051
rect 2881 218023 2909 218051
rect 2943 218023 2971 218051
rect 2757 217961 2785 217989
rect 2819 217961 2847 217989
rect 2881 217961 2909 217989
rect 2943 217961 2971 217989
rect 2757 209147 2785 209175
rect 2819 209147 2847 209175
rect 2881 209147 2909 209175
rect 2943 209147 2971 209175
rect 2757 209085 2785 209113
rect 2819 209085 2847 209113
rect 2881 209085 2909 209113
rect 2943 209085 2971 209113
rect 2757 209023 2785 209051
rect 2819 209023 2847 209051
rect 2881 209023 2909 209051
rect 2943 209023 2971 209051
rect 2757 208961 2785 208989
rect 2819 208961 2847 208989
rect 2881 208961 2909 208989
rect 2943 208961 2971 208989
rect 4617 299058 4645 299086
rect 4679 299058 4707 299086
rect 4741 299058 4769 299086
rect 4803 299058 4831 299086
rect 4617 298996 4645 299024
rect 4679 298996 4707 299024
rect 4741 298996 4769 299024
rect 4803 298996 4831 299024
rect 4617 298934 4645 298962
rect 4679 298934 4707 298962
rect 4741 298934 4769 298962
rect 4803 298934 4831 298962
rect 4617 298872 4645 298900
rect 4679 298872 4707 298900
rect 4741 298872 4769 298900
rect 4803 298872 4831 298900
rect 4617 293147 4645 293175
rect 4679 293147 4707 293175
rect 4741 293147 4769 293175
rect 4803 293147 4831 293175
rect 4617 293085 4645 293113
rect 4679 293085 4707 293113
rect 4741 293085 4769 293113
rect 4803 293085 4831 293113
rect 4617 293023 4645 293051
rect 4679 293023 4707 293051
rect 4741 293023 4769 293051
rect 4803 293023 4831 293051
rect 4617 292961 4645 292989
rect 4679 292961 4707 292989
rect 4741 292961 4769 292989
rect 4803 292961 4831 292989
rect 4617 284147 4645 284175
rect 4679 284147 4707 284175
rect 4741 284147 4769 284175
rect 4803 284147 4831 284175
rect 4617 284085 4645 284113
rect 4679 284085 4707 284113
rect 4741 284085 4769 284113
rect 4803 284085 4831 284113
rect 4617 284023 4645 284051
rect 4679 284023 4707 284051
rect 4741 284023 4769 284051
rect 4803 284023 4831 284051
rect 4617 283961 4645 283989
rect 4679 283961 4707 283989
rect 4741 283961 4769 283989
rect 4803 283961 4831 283989
rect 4617 275147 4645 275175
rect 4679 275147 4707 275175
rect 4741 275147 4769 275175
rect 4803 275147 4831 275175
rect 4617 275085 4645 275113
rect 4679 275085 4707 275113
rect 4741 275085 4769 275113
rect 4803 275085 4831 275113
rect 4617 275023 4645 275051
rect 4679 275023 4707 275051
rect 4741 275023 4769 275051
rect 4803 275023 4831 275051
rect 4617 274961 4645 274989
rect 4679 274961 4707 274989
rect 4741 274961 4769 274989
rect 4803 274961 4831 274989
rect 4617 266147 4645 266175
rect 4679 266147 4707 266175
rect 4741 266147 4769 266175
rect 4803 266147 4831 266175
rect 4617 266085 4645 266113
rect 4679 266085 4707 266113
rect 4741 266085 4769 266113
rect 4803 266085 4831 266113
rect 4617 266023 4645 266051
rect 4679 266023 4707 266051
rect 4741 266023 4769 266051
rect 4803 266023 4831 266051
rect 4617 265961 4645 265989
rect 4679 265961 4707 265989
rect 4741 265961 4769 265989
rect 4803 265961 4831 265989
rect 4617 257147 4645 257175
rect 4679 257147 4707 257175
rect 4741 257147 4769 257175
rect 4803 257147 4831 257175
rect 4617 257085 4645 257113
rect 4679 257085 4707 257113
rect 4741 257085 4769 257113
rect 4803 257085 4831 257113
rect 4617 257023 4645 257051
rect 4679 257023 4707 257051
rect 4741 257023 4769 257051
rect 4803 257023 4831 257051
rect 4617 256961 4645 256989
rect 4679 256961 4707 256989
rect 4741 256961 4769 256989
rect 4803 256961 4831 256989
rect 4617 248147 4645 248175
rect 4679 248147 4707 248175
rect 4741 248147 4769 248175
rect 4803 248147 4831 248175
rect 4617 248085 4645 248113
rect 4679 248085 4707 248113
rect 4741 248085 4769 248113
rect 4803 248085 4831 248113
rect 4617 248023 4645 248051
rect 4679 248023 4707 248051
rect 4741 248023 4769 248051
rect 4803 248023 4831 248051
rect 4617 247961 4645 247989
rect 4679 247961 4707 247989
rect 4741 247961 4769 247989
rect 4803 247961 4831 247989
rect 4617 239147 4645 239175
rect 4679 239147 4707 239175
rect 4741 239147 4769 239175
rect 4803 239147 4831 239175
rect 4617 239085 4645 239113
rect 4679 239085 4707 239113
rect 4741 239085 4769 239113
rect 4803 239085 4831 239113
rect 4617 239023 4645 239051
rect 4679 239023 4707 239051
rect 4741 239023 4769 239051
rect 4803 239023 4831 239051
rect 4617 238961 4645 238989
rect 4679 238961 4707 238989
rect 4741 238961 4769 238989
rect 4803 238961 4831 238989
rect 4617 230147 4645 230175
rect 4679 230147 4707 230175
rect 4741 230147 4769 230175
rect 4803 230147 4831 230175
rect 4617 230085 4645 230113
rect 4679 230085 4707 230113
rect 4741 230085 4769 230113
rect 4803 230085 4831 230113
rect 4617 230023 4645 230051
rect 4679 230023 4707 230051
rect 4741 230023 4769 230051
rect 4803 230023 4831 230051
rect 4617 229961 4645 229989
rect 4679 229961 4707 229989
rect 4741 229961 4769 229989
rect 4803 229961 4831 229989
rect 4617 221147 4645 221175
rect 4679 221147 4707 221175
rect 4741 221147 4769 221175
rect 4803 221147 4831 221175
rect 4617 221085 4645 221113
rect 4679 221085 4707 221113
rect 4741 221085 4769 221113
rect 4803 221085 4831 221113
rect 4617 221023 4645 221051
rect 4679 221023 4707 221051
rect 4741 221023 4769 221051
rect 4803 221023 4831 221051
rect 4617 220961 4645 220989
rect 4679 220961 4707 220989
rect 4741 220961 4769 220989
rect 4803 220961 4831 220989
rect 4617 212147 4645 212175
rect 4679 212147 4707 212175
rect 4741 212147 4769 212175
rect 4803 212147 4831 212175
rect 4617 212085 4645 212113
rect 4679 212085 4707 212113
rect 4741 212085 4769 212113
rect 4803 212085 4831 212113
rect 4617 212023 4645 212051
rect 4679 212023 4707 212051
rect 4741 212023 4769 212051
rect 4803 212023 4831 212051
rect 4617 211961 4645 211989
rect 4679 211961 4707 211989
rect 4741 211961 4769 211989
rect 4803 211961 4831 211989
rect 4617 203147 4645 203175
rect 4679 203147 4707 203175
rect 4741 203147 4769 203175
rect 4803 203147 4831 203175
rect 4617 203085 4645 203113
rect 4679 203085 4707 203113
rect 4741 203085 4769 203113
rect 4803 203085 4831 203113
rect 4617 203023 4645 203051
rect 4679 203023 4707 203051
rect 4741 203023 4769 203051
rect 4803 203023 4831 203051
rect 4617 202961 4645 202989
rect 4679 202961 4707 202989
rect 4741 202961 4769 202989
rect 4803 202961 4831 202989
rect 2757 200147 2785 200175
rect 2819 200147 2847 200175
rect 2881 200147 2909 200175
rect 2943 200147 2971 200175
rect 2757 200085 2785 200113
rect 2819 200085 2847 200113
rect 2881 200085 2909 200113
rect 2943 200085 2971 200113
rect 2757 200023 2785 200051
rect 2819 200023 2847 200051
rect 2881 200023 2909 200051
rect 2943 200023 2971 200051
rect 2757 199961 2785 199989
rect 2819 199961 2847 199989
rect 2881 199961 2909 199989
rect 2943 199961 2971 199989
rect 2757 191147 2785 191175
rect 2819 191147 2847 191175
rect 2881 191147 2909 191175
rect 2943 191147 2971 191175
rect 2757 191085 2785 191113
rect 2819 191085 2847 191113
rect 2881 191085 2909 191113
rect 2943 191085 2971 191113
rect 2757 191023 2785 191051
rect 2819 191023 2847 191051
rect 2881 191023 2909 191051
rect 2943 191023 2971 191051
rect 2757 190961 2785 190989
rect 2819 190961 2847 190989
rect 2881 190961 2909 190989
rect 2943 190961 2971 190989
rect 2757 182147 2785 182175
rect 2819 182147 2847 182175
rect 2881 182147 2909 182175
rect 2943 182147 2971 182175
rect 2757 182085 2785 182113
rect 2819 182085 2847 182113
rect 2881 182085 2909 182113
rect 2943 182085 2971 182113
rect 2757 182023 2785 182051
rect 2819 182023 2847 182051
rect 2881 182023 2909 182051
rect 2943 182023 2971 182051
rect 2757 181961 2785 181989
rect 2819 181961 2847 181989
rect 2881 181961 2909 181989
rect 2943 181961 2971 181989
rect -430 29147 -402 29175
rect -368 29147 -340 29175
rect -306 29147 -278 29175
rect -244 29147 -216 29175
rect -430 29085 -402 29113
rect -368 29085 -340 29113
rect -306 29085 -278 29113
rect -244 29085 -216 29113
rect -430 29023 -402 29051
rect -368 29023 -340 29051
rect -306 29023 -278 29051
rect -244 29023 -216 29051
rect -430 28961 -402 28989
rect -368 28961 -340 28989
rect -306 28961 -278 28989
rect -244 28961 -216 28989
rect -430 20147 -402 20175
rect -368 20147 -340 20175
rect -306 20147 -278 20175
rect -244 20147 -216 20175
rect -430 20085 -402 20113
rect -368 20085 -340 20113
rect -306 20085 -278 20113
rect -244 20085 -216 20113
rect -430 20023 -402 20051
rect -368 20023 -340 20051
rect -306 20023 -278 20051
rect -244 20023 -216 20051
rect -430 19961 -402 19989
rect -368 19961 -340 19989
rect -306 19961 -278 19989
rect -244 19961 -216 19989
rect 2757 173147 2785 173175
rect 2819 173147 2847 173175
rect 2881 173147 2909 173175
rect 2943 173147 2971 173175
rect 2757 173085 2785 173113
rect 2819 173085 2847 173113
rect 2881 173085 2909 173113
rect 2943 173085 2971 173113
rect 2757 173023 2785 173051
rect 2819 173023 2847 173051
rect 2881 173023 2909 173051
rect 2943 173023 2971 173051
rect 2757 172961 2785 172989
rect 2819 172961 2847 172989
rect 2881 172961 2909 172989
rect 2943 172961 2971 172989
rect 2757 164147 2785 164175
rect 2819 164147 2847 164175
rect 2881 164147 2909 164175
rect 2943 164147 2971 164175
rect 2757 164085 2785 164113
rect 2819 164085 2847 164113
rect 2881 164085 2909 164113
rect 2943 164085 2971 164113
rect 2757 164023 2785 164051
rect 2819 164023 2847 164051
rect 2881 164023 2909 164051
rect 2943 164023 2971 164051
rect 2757 163961 2785 163989
rect 2819 163961 2847 163989
rect 2881 163961 2909 163989
rect 2943 163961 2971 163989
rect 2757 155147 2785 155175
rect 2819 155147 2847 155175
rect 2881 155147 2909 155175
rect 2943 155147 2971 155175
rect 2757 155085 2785 155113
rect 2819 155085 2847 155113
rect 2881 155085 2909 155113
rect 2943 155085 2971 155113
rect 2757 155023 2785 155051
rect 2819 155023 2847 155051
rect 2881 155023 2909 155051
rect 2943 155023 2971 155051
rect 2757 154961 2785 154989
rect 2819 154961 2847 154989
rect 2881 154961 2909 154989
rect 2943 154961 2971 154989
rect 2757 146147 2785 146175
rect 2819 146147 2847 146175
rect 2881 146147 2909 146175
rect 2943 146147 2971 146175
rect 2757 146085 2785 146113
rect 2819 146085 2847 146113
rect 2881 146085 2909 146113
rect 2943 146085 2971 146113
rect 2757 146023 2785 146051
rect 2819 146023 2847 146051
rect 2881 146023 2909 146051
rect 2943 146023 2971 146051
rect 2757 145961 2785 145989
rect 2819 145961 2847 145989
rect 2881 145961 2909 145989
rect 2943 145961 2971 145989
rect 2757 137147 2785 137175
rect 2819 137147 2847 137175
rect 2881 137147 2909 137175
rect 2943 137147 2971 137175
rect 2757 137085 2785 137113
rect 2819 137085 2847 137113
rect 2881 137085 2909 137113
rect 2943 137085 2971 137113
rect 2757 137023 2785 137051
rect 2819 137023 2847 137051
rect 2881 137023 2909 137051
rect 2943 137023 2971 137051
rect 2757 136961 2785 136989
rect 2819 136961 2847 136989
rect 2881 136961 2909 136989
rect 2943 136961 2971 136989
rect 2757 128147 2785 128175
rect 2819 128147 2847 128175
rect 2881 128147 2909 128175
rect 2943 128147 2971 128175
rect 2757 128085 2785 128113
rect 2819 128085 2847 128113
rect 2881 128085 2909 128113
rect 2943 128085 2971 128113
rect 2757 128023 2785 128051
rect 2819 128023 2847 128051
rect 2881 128023 2909 128051
rect 2943 128023 2971 128051
rect 2757 127961 2785 127989
rect 2819 127961 2847 127989
rect 2881 127961 2909 127989
rect 2943 127961 2971 127989
rect 2757 119147 2785 119175
rect 2819 119147 2847 119175
rect 2881 119147 2909 119175
rect 2943 119147 2971 119175
rect 2757 119085 2785 119113
rect 2819 119085 2847 119113
rect 2881 119085 2909 119113
rect 2943 119085 2971 119113
rect 2757 119023 2785 119051
rect 2819 119023 2847 119051
rect 2881 119023 2909 119051
rect 2943 119023 2971 119051
rect 2757 118961 2785 118989
rect 2819 118961 2847 118989
rect 2881 118961 2909 118989
rect 2943 118961 2971 118989
rect 2757 110147 2785 110175
rect 2819 110147 2847 110175
rect 2881 110147 2909 110175
rect 2943 110147 2971 110175
rect 2757 110085 2785 110113
rect 2819 110085 2847 110113
rect 2881 110085 2909 110113
rect 2943 110085 2971 110113
rect 2757 110023 2785 110051
rect 2819 110023 2847 110051
rect 2881 110023 2909 110051
rect 2943 110023 2971 110051
rect 2757 109961 2785 109989
rect 2819 109961 2847 109989
rect 2881 109961 2909 109989
rect 2943 109961 2971 109989
rect -430 11147 -402 11175
rect -368 11147 -340 11175
rect -306 11147 -278 11175
rect -244 11147 -216 11175
rect -430 11085 -402 11113
rect -368 11085 -340 11113
rect -306 11085 -278 11113
rect -244 11085 -216 11113
rect -430 11023 -402 11051
rect -368 11023 -340 11051
rect -306 11023 -278 11051
rect -244 11023 -216 11051
rect -430 10961 -402 10989
rect -368 10961 -340 10989
rect -306 10961 -278 10989
rect -244 10961 -216 10989
rect 2757 101147 2785 101175
rect 2819 101147 2847 101175
rect 2881 101147 2909 101175
rect 2943 101147 2971 101175
rect 2757 101085 2785 101113
rect 2819 101085 2847 101113
rect 2881 101085 2909 101113
rect 2943 101085 2971 101113
rect 2757 101023 2785 101051
rect 2819 101023 2847 101051
rect 2881 101023 2909 101051
rect 2943 101023 2971 101051
rect 2757 100961 2785 100989
rect 2819 100961 2847 100989
rect 2881 100961 2909 100989
rect 2943 100961 2971 100989
rect 4617 194147 4645 194175
rect 4679 194147 4707 194175
rect 4741 194147 4769 194175
rect 4803 194147 4831 194175
rect 4617 194085 4645 194113
rect 4679 194085 4707 194113
rect 4741 194085 4769 194113
rect 4803 194085 4831 194113
rect 4617 194023 4645 194051
rect 4679 194023 4707 194051
rect 4741 194023 4769 194051
rect 4803 194023 4831 194051
rect 4617 193961 4645 193989
rect 4679 193961 4707 193989
rect 4741 193961 4769 193989
rect 4803 193961 4831 193989
rect 4617 185147 4645 185175
rect 4679 185147 4707 185175
rect 4741 185147 4769 185175
rect 4803 185147 4831 185175
rect 4617 185085 4645 185113
rect 4679 185085 4707 185113
rect 4741 185085 4769 185113
rect 4803 185085 4831 185113
rect 4617 185023 4645 185051
rect 4679 185023 4707 185051
rect 4741 185023 4769 185051
rect 4803 185023 4831 185051
rect 4617 184961 4645 184989
rect 4679 184961 4707 184989
rect 4741 184961 4769 184989
rect 4803 184961 4831 184989
rect 4617 176147 4645 176175
rect 4679 176147 4707 176175
rect 4741 176147 4769 176175
rect 4803 176147 4831 176175
rect 4617 176085 4645 176113
rect 4679 176085 4707 176113
rect 4741 176085 4769 176113
rect 4803 176085 4831 176113
rect 4617 176023 4645 176051
rect 4679 176023 4707 176051
rect 4741 176023 4769 176051
rect 4803 176023 4831 176051
rect 4617 175961 4645 175989
rect 4679 175961 4707 175989
rect 4741 175961 4769 175989
rect 4803 175961 4831 175989
rect 4617 167147 4645 167175
rect 4679 167147 4707 167175
rect 4741 167147 4769 167175
rect 4803 167147 4831 167175
rect 4617 167085 4645 167113
rect 4679 167085 4707 167113
rect 4741 167085 4769 167113
rect 4803 167085 4831 167113
rect 4617 167023 4645 167051
rect 4679 167023 4707 167051
rect 4741 167023 4769 167051
rect 4803 167023 4831 167051
rect 4617 166961 4645 166989
rect 4679 166961 4707 166989
rect 4741 166961 4769 166989
rect 4803 166961 4831 166989
rect 4617 158147 4645 158175
rect 4679 158147 4707 158175
rect 4741 158147 4769 158175
rect 4803 158147 4831 158175
rect 4617 158085 4645 158113
rect 4679 158085 4707 158113
rect 4741 158085 4769 158113
rect 4803 158085 4831 158113
rect 4617 158023 4645 158051
rect 4679 158023 4707 158051
rect 4741 158023 4769 158051
rect 4803 158023 4831 158051
rect 4617 157961 4645 157989
rect 4679 157961 4707 157989
rect 4741 157961 4769 157989
rect 4803 157961 4831 157989
rect 4617 149147 4645 149175
rect 4679 149147 4707 149175
rect 4741 149147 4769 149175
rect 4803 149147 4831 149175
rect 4617 149085 4645 149113
rect 4679 149085 4707 149113
rect 4741 149085 4769 149113
rect 4803 149085 4831 149113
rect 4617 149023 4645 149051
rect 4679 149023 4707 149051
rect 4741 149023 4769 149051
rect 4803 149023 4831 149051
rect 4617 148961 4645 148989
rect 4679 148961 4707 148989
rect 4741 148961 4769 148989
rect 4803 148961 4831 148989
rect 4617 140147 4645 140175
rect 4679 140147 4707 140175
rect 4741 140147 4769 140175
rect 4803 140147 4831 140175
rect 4617 140085 4645 140113
rect 4679 140085 4707 140113
rect 4741 140085 4769 140113
rect 4803 140085 4831 140113
rect 4617 140023 4645 140051
rect 4679 140023 4707 140051
rect 4741 140023 4769 140051
rect 4803 140023 4831 140051
rect 4617 139961 4645 139989
rect 4679 139961 4707 139989
rect 4741 139961 4769 139989
rect 4803 139961 4831 139989
rect 4617 131147 4645 131175
rect 4679 131147 4707 131175
rect 4741 131147 4769 131175
rect 4803 131147 4831 131175
rect 4617 131085 4645 131113
rect 4679 131085 4707 131113
rect 4741 131085 4769 131113
rect 4803 131085 4831 131113
rect 4617 131023 4645 131051
rect 4679 131023 4707 131051
rect 4741 131023 4769 131051
rect 4803 131023 4831 131051
rect 4617 130961 4645 130989
rect 4679 130961 4707 130989
rect 4741 130961 4769 130989
rect 4803 130961 4831 130989
rect 4617 122147 4645 122175
rect 4679 122147 4707 122175
rect 4741 122147 4769 122175
rect 4803 122147 4831 122175
rect 4617 122085 4645 122113
rect 4679 122085 4707 122113
rect 4741 122085 4769 122113
rect 4803 122085 4831 122113
rect 4617 122023 4645 122051
rect 4679 122023 4707 122051
rect 4741 122023 4769 122051
rect 4803 122023 4831 122051
rect 4617 121961 4645 121989
rect 4679 121961 4707 121989
rect 4741 121961 4769 121989
rect 4803 121961 4831 121989
rect 4617 113147 4645 113175
rect 4679 113147 4707 113175
rect 4741 113147 4769 113175
rect 4803 113147 4831 113175
rect 4617 113085 4645 113113
rect 4679 113085 4707 113113
rect 4741 113085 4769 113113
rect 4803 113085 4831 113113
rect 4617 113023 4645 113051
rect 4679 113023 4707 113051
rect 4741 113023 4769 113051
rect 4803 113023 4831 113051
rect 4617 112961 4645 112989
rect 4679 112961 4707 112989
rect 4741 112961 4769 112989
rect 4803 112961 4831 112989
rect 4617 104147 4645 104175
rect 4679 104147 4707 104175
rect 4741 104147 4769 104175
rect 4803 104147 4831 104175
rect 4617 104085 4645 104113
rect 4679 104085 4707 104113
rect 4741 104085 4769 104113
rect 4803 104085 4831 104113
rect 4617 104023 4645 104051
rect 4679 104023 4707 104051
rect 4741 104023 4769 104051
rect 4803 104023 4831 104051
rect 4617 103961 4645 103989
rect 4679 103961 4707 103989
rect 4741 103961 4769 103989
rect 4803 103961 4831 103989
rect 2757 92147 2785 92175
rect 2819 92147 2847 92175
rect 2881 92147 2909 92175
rect 2943 92147 2971 92175
rect 2757 92085 2785 92113
rect 2819 92085 2847 92113
rect 2881 92085 2909 92113
rect 2943 92085 2971 92113
rect 2757 92023 2785 92051
rect 2819 92023 2847 92051
rect 2881 92023 2909 92051
rect 2943 92023 2971 92051
rect 2757 91961 2785 91989
rect 2819 91961 2847 91989
rect 2881 91961 2909 91989
rect 2943 91961 2971 91989
rect 2757 83147 2785 83175
rect 2819 83147 2847 83175
rect 2881 83147 2909 83175
rect 2943 83147 2971 83175
rect 2757 83085 2785 83113
rect 2819 83085 2847 83113
rect 2881 83085 2909 83113
rect 2943 83085 2971 83113
rect 2757 83023 2785 83051
rect 2819 83023 2847 83051
rect 2881 83023 2909 83051
rect 2943 83023 2971 83051
rect 2757 82961 2785 82989
rect 2819 82961 2847 82989
rect 2881 82961 2909 82989
rect 2943 82961 2971 82989
rect 2757 74147 2785 74175
rect 2819 74147 2847 74175
rect 2881 74147 2909 74175
rect 2943 74147 2971 74175
rect 2757 74085 2785 74113
rect 2819 74085 2847 74113
rect 2881 74085 2909 74113
rect 2943 74085 2971 74113
rect 2757 74023 2785 74051
rect 2819 74023 2847 74051
rect 2881 74023 2909 74051
rect 2943 74023 2971 74051
rect 2757 73961 2785 73989
rect 2819 73961 2847 73989
rect 2881 73961 2909 73989
rect 2943 73961 2971 73989
rect 2757 65147 2785 65175
rect 2819 65147 2847 65175
rect 2881 65147 2909 65175
rect 2943 65147 2971 65175
rect 2757 65085 2785 65113
rect 2819 65085 2847 65113
rect 2881 65085 2909 65113
rect 2943 65085 2971 65113
rect 2757 65023 2785 65051
rect 2819 65023 2847 65051
rect 2881 65023 2909 65051
rect 2943 65023 2971 65051
rect 2757 64961 2785 64989
rect 2819 64961 2847 64989
rect 2881 64961 2909 64989
rect 2943 64961 2971 64989
rect 2757 56147 2785 56175
rect 2819 56147 2847 56175
rect 2881 56147 2909 56175
rect 2943 56147 2971 56175
rect 2757 56085 2785 56113
rect 2819 56085 2847 56113
rect 2881 56085 2909 56113
rect 2943 56085 2971 56113
rect 2757 56023 2785 56051
rect 2819 56023 2847 56051
rect 2881 56023 2909 56051
rect 2943 56023 2971 56051
rect 2757 55961 2785 55989
rect 2819 55961 2847 55989
rect 2881 55961 2909 55989
rect 2943 55961 2971 55989
rect 2757 47147 2785 47175
rect 2819 47147 2847 47175
rect 2881 47147 2909 47175
rect 2943 47147 2971 47175
rect 2757 47085 2785 47113
rect 2819 47085 2847 47113
rect 2881 47085 2909 47113
rect 2943 47085 2971 47113
rect 2757 47023 2785 47051
rect 2819 47023 2847 47051
rect 2881 47023 2909 47051
rect 2943 47023 2971 47051
rect 2757 46961 2785 46989
rect 2819 46961 2847 46989
rect 2881 46961 2909 46989
rect 2943 46961 2971 46989
rect 2757 38147 2785 38175
rect 2819 38147 2847 38175
rect 2881 38147 2909 38175
rect 2943 38147 2971 38175
rect 2757 38085 2785 38113
rect 2819 38085 2847 38113
rect 2881 38085 2909 38113
rect 2943 38085 2971 38113
rect 2757 38023 2785 38051
rect 2819 38023 2847 38051
rect 2881 38023 2909 38051
rect 2943 38023 2971 38051
rect 2757 37961 2785 37989
rect 2819 37961 2847 37989
rect 2881 37961 2909 37989
rect 2943 37961 2971 37989
rect 2757 29147 2785 29175
rect 2819 29147 2847 29175
rect 2881 29147 2909 29175
rect 2943 29147 2971 29175
rect 2757 29085 2785 29113
rect 2819 29085 2847 29113
rect 2881 29085 2909 29113
rect 2943 29085 2971 29113
rect 2757 29023 2785 29051
rect 2819 29023 2847 29051
rect 2881 29023 2909 29051
rect 2943 29023 2971 29051
rect 2757 28961 2785 28989
rect 2819 28961 2847 28989
rect 2881 28961 2909 28989
rect 2943 28961 2971 28989
rect 2757 20147 2785 20175
rect 2819 20147 2847 20175
rect 2881 20147 2909 20175
rect 2943 20147 2971 20175
rect 2757 20085 2785 20113
rect 2819 20085 2847 20113
rect 2881 20085 2909 20113
rect 2943 20085 2971 20113
rect 2757 20023 2785 20051
rect 2819 20023 2847 20051
rect 2881 20023 2909 20051
rect 2943 20023 2971 20051
rect 2757 19961 2785 19989
rect 2819 19961 2847 19989
rect 2881 19961 2909 19989
rect 2943 19961 2971 19989
rect 2757 11147 2785 11175
rect 2819 11147 2847 11175
rect 2881 11147 2909 11175
rect 2943 11147 2971 11175
rect 2757 11085 2785 11113
rect 2819 11085 2847 11113
rect 2881 11085 2909 11113
rect 2943 11085 2971 11113
rect 2757 11023 2785 11051
rect 2819 11023 2847 11051
rect 2881 11023 2909 11051
rect 2943 11023 2971 11051
rect 2757 10961 2785 10989
rect 2819 10961 2847 10989
rect 2881 10961 2909 10989
rect 2943 10961 2971 10989
rect -430 2147 -402 2175
rect -368 2147 -340 2175
rect -306 2147 -278 2175
rect -244 2147 -216 2175
rect -430 2085 -402 2113
rect -368 2085 -340 2113
rect -306 2085 -278 2113
rect -244 2085 -216 2113
rect -430 2023 -402 2051
rect -368 2023 -340 2051
rect -306 2023 -278 2051
rect -244 2023 -216 2051
rect -430 1961 -402 1989
rect -368 1961 -340 1989
rect -306 1961 -278 1989
rect -244 1961 -216 1989
rect -430 -108 -402 -80
rect -368 -108 -340 -80
rect -306 -108 -278 -80
rect -244 -108 -216 -80
rect -430 -170 -402 -142
rect -368 -170 -340 -142
rect -306 -170 -278 -142
rect -244 -170 -216 -142
rect -430 -232 -402 -204
rect -368 -232 -340 -204
rect -306 -232 -278 -204
rect -244 -232 -216 -204
rect -430 -294 -402 -266
rect -368 -294 -340 -266
rect -306 -294 -278 -266
rect -244 -294 -216 -266
rect 2757 2147 2785 2175
rect 2819 2147 2847 2175
rect 2881 2147 2909 2175
rect 2943 2147 2971 2175
rect 2757 2085 2785 2113
rect 2819 2085 2847 2113
rect 2881 2085 2909 2113
rect 2943 2085 2971 2113
rect 2757 2023 2785 2051
rect 2819 2023 2847 2051
rect 2881 2023 2909 2051
rect 2943 2023 2971 2051
rect 2757 1961 2785 1989
rect 2819 1961 2847 1989
rect 2881 1961 2909 1989
rect 2943 1961 2971 1989
rect 2757 -108 2785 -80
rect 2819 -108 2847 -80
rect 2881 -108 2909 -80
rect 2943 -108 2971 -80
rect 2757 -170 2785 -142
rect 2819 -170 2847 -142
rect 2881 -170 2909 -142
rect 2943 -170 2971 -142
rect 2757 -232 2785 -204
rect 2819 -232 2847 -204
rect 2881 -232 2909 -204
rect 2943 -232 2971 -204
rect 2757 -294 2785 -266
rect 2819 -294 2847 -266
rect 2881 -294 2909 -266
rect 2943 -294 2971 -266
rect -910 -588 -882 -560
rect -848 -588 -820 -560
rect -786 -588 -758 -560
rect -724 -588 -696 -560
rect -910 -650 -882 -622
rect -848 -650 -820 -622
rect -786 -650 -758 -622
rect -724 -650 -696 -622
rect -910 -712 -882 -684
rect -848 -712 -820 -684
rect -786 -712 -758 -684
rect -724 -712 -696 -684
rect -910 -774 -882 -746
rect -848 -774 -820 -746
rect -786 -774 -758 -746
rect -724 -774 -696 -746
rect 4617 95147 4645 95175
rect 4679 95147 4707 95175
rect 4741 95147 4769 95175
rect 4803 95147 4831 95175
rect 4617 95085 4645 95113
rect 4679 95085 4707 95113
rect 4741 95085 4769 95113
rect 4803 95085 4831 95113
rect 4617 95023 4645 95051
rect 4679 95023 4707 95051
rect 4741 95023 4769 95051
rect 4803 95023 4831 95051
rect 4617 94961 4645 94989
rect 4679 94961 4707 94989
rect 4741 94961 4769 94989
rect 4803 94961 4831 94989
rect 4617 86147 4645 86175
rect 4679 86147 4707 86175
rect 4741 86147 4769 86175
rect 4803 86147 4831 86175
rect 4617 86085 4645 86113
rect 4679 86085 4707 86113
rect 4741 86085 4769 86113
rect 4803 86085 4831 86113
rect 4617 86023 4645 86051
rect 4679 86023 4707 86051
rect 4741 86023 4769 86051
rect 4803 86023 4831 86051
rect 4617 85961 4645 85989
rect 4679 85961 4707 85989
rect 4741 85961 4769 85989
rect 4803 85961 4831 85989
rect 4617 77147 4645 77175
rect 4679 77147 4707 77175
rect 4741 77147 4769 77175
rect 4803 77147 4831 77175
rect 4617 77085 4645 77113
rect 4679 77085 4707 77113
rect 4741 77085 4769 77113
rect 4803 77085 4831 77113
rect 4617 77023 4645 77051
rect 4679 77023 4707 77051
rect 4741 77023 4769 77051
rect 4803 77023 4831 77051
rect 4617 76961 4645 76989
rect 4679 76961 4707 76989
rect 4741 76961 4769 76989
rect 4803 76961 4831 76989
rect 4617 68147 4645 68175
rect 4679 68147 4707 68175
rect 4741 68147 4769 68175
rect 4803 68147 4831 68175
rect 4617 68085 4645 68113
rect 4679 68085 4707 68113
rect 4741 68085 4769 68113
rect 4803 68085 4831 68113
rect 4617 68023 4645 68051
rect 4679 68023 4707 68051
rect 4741 68023 4769 68051
rect 4803 68023 4831 68051
rect 4617 67961 4645 67989
rect 4679 67961 4707 67989
rect 4741 67961 4769 67989
rect 4803 67961 4831 67989
rect 4617 59147 4645 59175
rect 4679 59147 4707 59175
rect 4741 59147 4769 59175
rect 4803 59147 4831 59175
rect 4617 59085 4645 59113
rect 4679 59085 4707 59113
rect 4741 59085 4769 59113
rect 4803 59085 4831 59113
rect 4617 59023 4645 59051
rect 4679 59023 4707 59051
rect 4741 59023 4769 59051
rect 4803 59023 4831 59051
rect 4617 58961 4645 58989
rect 4679 58961 4707 58989
rect 4741 58961 4769 58989
rect 4803 58961 4831 58989
rect 4617 50147 4645 50175
rect 4679 50147 4707 50175
rect 4741 50147 4769 50175
rect 4803 50147 4831 50175
rect 4617 50085 4645 50113
rect 4679 50085 4707 50113
rect 4741 50085 4769 50113
rect 4803 50085 4831 50113
rect 4617 50023 4645 50051
rect 4679 50023 4707 50051
rect 4741 50023 4769 50051
rect 4803 50023 4831 50051
rect 4617 49961 4645 49989
rect 4679 49961 4707 49989
rect 4741 49961 4769 49989
rect 4803 49961 4831 49989
rect 4617 41147 4645 41175
rect 4679 41147 4707 41175
rect 4741 41147 4769 41175
rect 4803 41147 4831 41175
rect 4617 41085 4645 41113
rect 4679 41085 4707 41113
rect 4741 41085 4769 41113
rect 4803 41085 4831 41113
rect 4617 41023 4645 41051
rect 4679 41023 4707 41051
rect 4741 41023 4769 41051
rect 4803 41023 4831 41051
rect 4617 40961 4645 40989
rect 4679 40961 4707 40989
rect 4741 40961 4769 40989
rect 4803 40961 4831 40989
rect 4617 32147 4645 32175
rect 4679 32147 4707 32175
rect 4741 32147 4769 32175
rect 4803 32147 4831 32175
rect 4617 32085 4645 32113
rect 4679 32085 4707 32113
rect 4741 32085 4769 32113
rect 4803 32085 4831 32113
rect 4617 32023 4645 32051
rect 4679 32023 4707 32051
rect 4741 32023 4769 32051
rect 4803 32023 4831 32051
rect 4617 31961 4645 31989
rect 4679 31961 4707 31989
rect 4741 31961 4769 31989
rect 4803 31961 4831 31989
rect 4617 23147 4645 23175
rect 4679 23147 4707 23175
rect 4741 23147 4769 23175
rect 4803 23147 4831 23175
rect 4617 23085 4645 23113
rect 4679 23085 4707 23113
rect 4741 23085 4769 23113
rect 4803 23085 4831 23113
rect 4617 23023 4645 23051
rect 4679 23023 4707 23051
rect 4741 23023 4769 23051
rect 4803 23023 4831 23051
rect 4617 22961 4645 22989
rect 4679 22961 4707 22989
rect 4741 22961 4769 22989
rect 4803 22961 4831 22989
rect 4617 14147 4645 14175
rect 4679 14147 4707 14175
rect 4741 14147 4769 14175
rect 4803 14147 4831 14175
rect 4617 14085 4645 14113
rect 4679 14085 4707 14113
rect 4741 14085 4769 14113
rect 4803 14085 4831 14113
rect 4617 14023 4645 14051
rect 4679 14023 4707 14051
rect 4741 14023 4769 14051
rect 4803 14023 4831 14051
rect 4617 13961 4645 13989
rect 4679 13961 4707 13989
rect 4741 13961 4769 13989
rect 4803 13961 4831 13989
rect 4617 5147 4645 5175
rect 4679 5147 4707 5175
rect 4741 5147 4769 5175
rect 4803 5147 4831 5175
rect 4617 5085 4645 5113
rect 4679 5085 4707 5113
rect 4741 5085 4769 5113
rect 4803 5085 4831 5113
rect 4617 5023 4645 5051
rect 4679 5023 4707 5051
rect 4741 5023 4769 5051
rect 4803 5023 4831 5051
rect 4617 4961 4645 4989
rect 4679 4961 4707 4989
rect 4741 4961 4769 4989
rect 4803 4961 4831 4989
rect 4617 -588 4645 -560
rect 4679 -588 4707 -560
rect 4741 -588 4769 -560
rect 4803 -588 4831 -560
rect 4617 -650 4645 -622
rect 4679 -650 4707 -622
rect 4741 -650 4769 -622
rect 4803 -650 4831 -622
rect 4617 -712 4645 -684
rect 4679 -712 4707 -684
rect 4741 -712 4769 -684
rect 4803 -712 4831 -684
rect 4617 -774 4645 -746
rect 4679 -774 4707 -746
rect 4741 -774 4769 -746
rect 4803 -774 4831 -746
rect 18117 298578 18145 298606
rect 18179 298578 18207 298606
rect 18241 298578 18269 298606
rect 18303 298578 18331 298606
rect 18117 298516 18145 298544
rect 18179 298516 18207 298544
rect 18241 298516 18269 298544
rect 18303 298516 18331 298544
rect 18117 298454 18145 298482
rect 18179 298454 18207 298482
rect 18241 298454 18269 298482
rect 18303 298454 18331 298482
rect 18117 298392 18145 298420
rect 18179 298392 18207 298420
rect 18241 298392 18269 298420
rect 18303 298392 18331 298420
rect 18117 290147 18145 290175
rect 18179 290147 18207 290175
rect 18241 290147 18269 290175
rect 18303 290147 18331 290175
rect 18117 290085 18145 290113
rect 18179 290085 18207 290113
rect 18241 290085 18269 290113
rect 18303 290085 18331 290113
rect 18117 290023 18145 290051
rect 18179 290023 18207 290051
rect 18241 290023 18269 290051
rect 18303 290023 18331 290051
rect 18117 289961 18145 289989
rect 18179 289961 18207 289989
rect 18241 289961 18269 289989
rect 18303 289961 18331 289989
rect 18117 281147 18145 281175
rect 18179 281147 18207 281175
rect 18241 281147 18269 281175
rect 18303 281147 18331 281175
rect 18117 281085 18145 281113
rect 18179 281085 18207 281113
rect 18241 281085 18269 281113
rect 18303 281085 18331 281113
rect 18117 281023 18145 281051
rect 18179 281023 18207 281051
rect 18241 281023 18269 281051
rect 18303 281023 18331 281051
rect 18117 280961 18145 280989
rect 18179 280961 18207 280989
rect 18241 280961 18269 280989
rect 18303 280961 18331 280989
rect 18117 272147 18145 272175
rect 18179 272147 18207 272175
rect 18241 272147 18269 272175
rect 18303 272147 18331 272175
rect 18117 272085 18145 272113
rect 18179 272085 18207 272113
rect 18241 272085 18269 272113
rect 18303 272085 18331 272113
rect 18117 272023 18145 272051
rect 18179 272023 18207 272051
rect 18241 272023 18269 272051
rect 18303 272023 18331 272051
rect 18117 271961 18145 271989
rect 18179 271961 18207 271989
rect 18241 271961 18269 271989
rect 18303 271961 18331 271989
rect 18117 263147 18145 263175
rect 18179 263147 18207 263175
rect 18241 263147 18269 263175
rect 18303 263147 18331 263175
rect 18117 263085 18145 263113
rect 18179 263085 18207 263113
rect 18241 263085 18269 263113
rect 18303 263085 18331 263113
rect 18117 263023 18145 263051
rect 18179 263023 18207 263051
rect 18241 263023 18269 263051
rect 18303 263023 18331 263051
rect 18117 262961 18145 262989
rect 18179 262961 18207 262989
rect 18241 262961 18269 262989
rect 18303 262961 18331 262989
rect 18117 254147 18145 254175
rect 18179 254147 18207 254175
rect 18241 254147 18269 254175
rect 18303 254147 18331 254175
rect 18117 254085 18145 254113
rect 18179 254085 18207 254113
rect 18241 254085 18269 254113
rect 18303 254085 18331 254113
rect 18117 254023 18145 254051
rect 18179 254023 18207 254051
rect 18241 254023 18269 254051
rect 18303 254023 18331 254051
rect 18117 253961 18145 253989
rect 18179 253961 18207 253989
rect 18241 253961 18269 253989
rect 18303 253961 18331 253989
rect 18117 245147 18145 245175
rect 18179 245147 18207 245175
rect 18241 245147 18269 245175
rect 18303 245147 18331 245175
rect 18117 245085 18145 245113
rect 18179 245085 18207 245113
rect 18241 245085 18269 245113
rect 18303 245085 18331 245113
rect 18117 245023 18145 245051
rect 18179 245023 18207 245051
rect 18241 245023 18269 245051
rect 18303 245023 18331 245051
rect 18117 244961 18145 244989
rect 18179 244961 18207 244989
rect 18241 244961 18269 244989
rect 18303 244961 18331 244989
rect 18117 236147 18145 236175
rect 18179 236147 18207 236175
rect 18241 236147 18269 236175
rect 18303 236147 18331 236175
rect 18117 236085 18145 236113
rect 18179 236085 18207 236113
rect 18241 236085 18269 236113
rect 18303 236085 18331 236113
rect 18117 236023 18145 236051
rect 18179 236023 18207 236051
rect 18241 236023 18269 236051
rect 18303 236023 18331 236051
rect 18117 235961 18145 235989
rect 18179 235961 18207 235989
rect 18241 235961 18269 235989
rect 18303 235961 18331 235989
rect 18117 227147 18145 227175
rect 18179 227147 18207 227175
rect 18241 227147 18269 227175
rect 18303 227147 18331 227175
rect 18117 227085 18145 227113
rect 18179 227085 18207 227113
rect 18241 227085 18269 227113
rect 18303 227085 18331 227113
rect 18117 227023 18145 227051
rect 18179 227023 18207 227051
rect 18241 227023 18269 227051
rect 18303 227023 18331 227051
rect 18117 226961 18145 226989
rect 18179 226961 18207 226989
rect 18241 226961 18269 226989
rect 18303 226961 18331 226989
rect 18117 218147 18145 218175
rect 18179 218147 18207 218175
rect 18241 218147 18269 218175
rect 18303 218147 18331 218175
rect 18117 218085 18145 218113
rect 18179 218085 18207 218113
rect 18241 218085 18269 218113
rect 18303 218085 18331 218113
rect 18117 218023 18145 218051
rect 18179 218023 18207 218051
rect 18241 218023 18269 218051
rect 18303 218023 18331 218051
rect 18117 217961 18145 217989
rect 18179 217961 18207 217989
rect 18241 217961 18269 217989
rect 18303 217961 18331 217989
rect 18117 209147 18145 209175
rect 18179 209147 18207 209175
rect 18241 209147 18269 209175
rect 18303 209147 18331 209175
rect 18117 209085 18145 209113
rect 18179 209085 18207 209113
rect 18241 209085 18269 209113
rect 18303 209085 18331 209113
rect 18117 209023 18145 209051
rect 18179 209023 18207 209051
rect 18241 209023 18269 209051
rect 18303 209023 18331 209051
rect 18117 208961 18145 208989
rect 18179 208961 18207 208989
rect 18241 208961 18269 208989
rect 18303 208961 18331 208989
rect 18117 200147 18145 200175
rect 18179 200147 18207 200175
rect 18241 200147 18269 200175
rect 18303 200147 18331 200175
rect 18117 200085 18145 200113
rect 18179 200085 18207 200113
rect 18241 200085 18269 200113
rect 18303 200085 18331 200113
rect 18117 200023 18145 200051
rect 18179 200023 18207 200051
rect 18241 200023 18269 200051
rect 18303 200023 18331 200051
rect 18117 199961 18145 199989
rect 18179 199961 18207 199989
rect 18241 199961 18269 199989
rect 18303 199961 18331 199989
rect 18117 191147 18145 191175
rect 18179 191147 18207 191175
rect 18241 191147 18269 191175
rect 18303 191147 18331 191175
rect 18117 191085 18145 191113
rect 18179 191085 18207 191113
rect 18241 191085 18269 191113
rect 18303 191085 18331 191113
rect 18117 191023 18145 191051
rect 18179 191023 18207 191051
rect 18241 191023 18269 191051
rect 18303 191023 18331 191051
rect 18117 190961 18145 190989
rect 18179 190961 18207 190989
rect 18241 190961 18269 190989
rect 18303 190961 18331 190989
rect 18117 182147 18145 182175
rect 18179 182147 18207 182175
rect 18241 182147 18269 182175
rect 18303 182147 18331 182175
rect 18117 182085 18145 182113
rect 18179 182085 18207 182113
rect 18241 182085 18269 182113
rect 18303 182085 18331 182113
rect 18117 182023 18145 182051
rect 18179 182023 18207 182051
rect 18241 182023 18269 182051
rect 18303 182023 18331 182051
rect 18117 181961 18145 181989
rect 18179 181961 18207 181989
rect 18241 181961 18269 181989
rect 18303 181961 18331 181989
rect 18117 173147 18145 173175
rect 18179 173147 18207 173175
rect 18241 173147 18269 173175
rect 18303 173147 18331 173175
rect 18117 173085 18145 173113
rect 18179 173085 18207 173113
rect 18241 173085 18269 173113
rect 18303 173085 18331 173113
rect 18117 173023 18145 173051
rect 18179 173023 18207 173051
rect 18241 173023 18269 173051
rect 18303 173023 18331 173051
rect 18117 172961 18145 172989
rect 18179 172961 18207 172989
rect 18241 172961 18269 172989
rect 18303 172961 18331 172989
rect 18117 164147 18145 164175
rect 18179 164147 18207 164175
rect 18241 164147 18269 164175
rect 18303 164147 18331 164175
rect 18117 164085 18145 164113
rect 18179 164085 18207 164113
rect 18241 164085 18269 164113
rect 18303 164085 18331 164113
rect 18117 164023 18145 164051
rect 18179 164023 18207 164051
rect 18241 164023 18269 164051
rect 18303 164023 18331 164051
rect 18117 163961 18145 163989
rect 18179 163961 18207 163989
rect 18241 163961 18269 163989
rect 18303 163961 18331 163989
rect 18117 155147 18145 155175
rect 18179 155147 18207 155175
rect 18241 155147 18269 155175
rect 18303 155147 18331 155175
rect 18117 155085 18145 155113
rect 18179 155085 18207 155113
rect 18241 155085 18269 155113
rect 18303 155085 18331 155113
rect 18117 155023 18145 155051
rect 18179 155023 18207 155051
rect 18241 155023 18269 155051
rect 18303 155023 18331 155051
rect 18117 154961 18145 154989
rect 18179 154961 18207 154989
rect 18241 154961 18269 154989
rect 18303 154961 18331 154989
rect 18117 146147 18145 146175
rect 18179 146147 18207 146175
rect 18241 146147 18269 146175
rect 18303 146147 18331 146175
rect 18117 146085 18145 146113
rect 18179 146085 18207 146113
rect 18241 146085 18269 146113
rect 18303 146085 18331 146113
rect 18117 146023 18145 146051
rect 18179 146023 18207 146051
rect 18241 146023 18269 146051
rect 18303 146023 18331 146051
rect 18117 145961 18145 145989
rect 18179 145961 18207 145989
rect 18241 145961 18269 145989
rect 18303 145961 18331 145989
rect 18117 137147 18145 137175
rect 18179 137147 18207 137175
rect 18241 137147 18269 137175
rect 18303 137147 18331 137175
rect 18117 137085 18145 137113
rect 18179 137085 18207 137113
rect 18241 137085 18269 137113
rect 18303 137085 18331 137113
rect 18117 137023 18145 137051
rect 18179 137023 18207 137051
rect 18241 137023 18269 137051
rect 18303 137023 18331 137051
rect 18117 136961 18145 136989
rect 18179 136961 18207 136989
rect 18241 136961 18269 136989
rect 18303 136961 18331 136989
rect 18117 128147 18145 128175
rect 18179 128147 18207 128175
rect 18241 128147 18269 128175
rect 18303 128147 18331 128175
rect 18117 128085 18145 128113
rect 18179 128085 18207 128113
rect 18241 128085 18269 128113
rect 18303 128085 18331 128113
rect 18117 128023 18145 128051
rect 18179 128023 18207 128051
rect 18241 128023 18269 128051
rect 18303 128023 18331 128051
rect 18117 127961 18145 127989
rect 18179 127961 18207 127989
rect 18241 127961 18269 127989
rect 18303 127961 18331 127989
rect 18117 119147 18145 119175
rect 18179 119147 18207 119175
rect 18241 119147 18269 119175
rect 18303 119147 18331 119175
rect 18117 119085 18145 119113
rect 18179 119085 18207 119113
rect 18241 119085 18269 119113
rect 18303 119085 18331 119113
rect 18117 119023 18145 119051
rect 18179 119023 18207 119051
rect 18241 119023 18269 119051
rect 18303 119023 18331 119051
rect 18117 118961 18145 118989
rect 18179 118961 18207 118989
rect 18241 118961 18269 118989
rect 18303 118961 18331 118989
rect 18117 110147 18145 110175
rect 18179 110147 18207 110175
rect 18241 110147 18269 110175
rect 18303 110147 18331 110175
rect 18117 110085 18145 110113
rect 18179 110085 18207 110113
rect 18241 110085 18269 110113
rect 18303 110085 18331 110113
rect 18117 110023 18145 110051
rect 18179 110023 18207 110051
rect 18241 110023 18269 110051
rect 18303 110023 18331 110051
rect 18117 109961 18145 109989
rect 18179 109961 18207 109989
rect 18241 109961 18269 109989
rect 18303 109961 18331 109989
rect 18117 101147 18145 101175
rect 18179 101147 18207 101175
rect 18241 101147 18269 101175
rect 18303 101147 18331 101175
rect 18117 101085 18145 101113
rect 18179 101085 18207 101113
rect 18241 101085 18269 101113
rect 18303 101085 18331 101113
rect 18117 101023 18145 101051
rect 18179 101023 18207 101051
rect 18241 101023 18269 101051
rect 18303 101023 18331 101051
rect 18117 100961 18145 100989
rect 18179 100961 18207 100989
rect 18241 100961 18269 100989
rect 18303 100961 18331 100989
rect 18117 92147 18145 92175
rect 18179 92147 18207 92175
rect 18241 92147 18269 92175
rect 18303 92147 18331 92175
rect 18117 92085 18145 92113
rect 18179 92085 18207 92113
rect 18241 92085 18269 92113
rect 18303 92085 18331 92113
rect 18117 92023 18145 92051
rect 18179 92023 18207 92051
rect 18241 92023 18269 92051
rect 18303 92023 18331 92051
rect 18117 91961 18145 91989
rect 18179 91961 18207 91989
rect 18241 91961 18269 91989
rect 18303 91961 18331 91989
rect 18117 83147 18145 83175
rect 18179 83147 18207 83175
rect 18241 83147 18269 83175
rect 18303 83147 18331 83175
rect 18117 83085 18145 83113
rect 18179 83085 18207 83113
rect 18241 83085 18269 83113
rect 18303 83085 18331 83113
rect 18117 83023 18145 83051
rect 18179 83023 18207 83051
rect 18241 83023 18269 83051
rect 18303 83023 18331 83051
rect 18117 82961 18145 82989
rect 18179 82961 18207 82989
rect 18241 82961 18269 82989
rect 18303 82961 18331 82989
rect 18117 74147 18145 74175
rect 18179 74147 18207 74175
rect 18241 74147 18269 74175
rect 18303 74147 18331 74175
rect 18117 74085 18145 74113
rect 18179 74085 18207 74113
rect 18241 74085 18269 74113
rect 18303 74085 18331 74113
rect 18117 74023 18145 74051
rect 18179 74023 18207 74051
rect 18241 74023 18269 74051
rect 18303 74023 18331 74051
rect 18117 73961 18145 73989
rect 18179 73961 18207 73989
rect 18241 73961 18269 73989
rect 18303 73961 18331 73989
rect 18117 65147 18145 65175
rect 18179 65147 18207 65175
rect 18241 65147 18269 65175
rect 18303 65147 18331 65175
rect 18117 65085 18145 65113
rect 18179 65085 18207 65113
rect 18241 65085 18269 65113
rect 18303 65085 18331 65113
rect 18117 65023 18145 65051
rect 18179 65023 18207 65051
rect 18241 65023 18269 65051
rect 18303 65023 18331 65051
rect 18117 64961 18145 64989
rect 18179 64961 18207 64989
rect 18241 64961 18269 64989
rect 18303 64961 18331 64989
rect 18117 56147 18145 56175
rect 18179 56147 18207 56175
rect 18241 56147 18269 56175
rect 18303 56147 18331 56175
rect 18117 56085 18145 56113
rect 18179 56085 18207 56113
rect 18241 56085 18269 56113
rect 18303 56085 18331 56113
rect 18117 56023 18145 56051
rect 18179 56023 18207 56051
rect 18241 56023 18269 56051
rect 18303 56023 18331 56051
rect 18117 55961 18145 55989
rect 18179 55961 18207 55989
rect 18241 55961 18269 55989
rect 18303 55961 18331 55989
rect 18117 47147 18145 47175
rect 18179 47147 18207 47175
rect 18241 47147 18269 47175
rect 18303 47147 18331 47175
rect 18117 47085 18145 47113
rect 18179 47085 18207 47113
rect 18241 47085 18269 47113
rect 18303 47085 18331 47113
rect 18117 47023 18145 47051
rect 18179 47023 18207 47051
rect 18241 47023 18269 47051
rect 18303 47023 18331 47051
rect 18117 46961 18145 46989
rect 18179 46961 18207 46989
rect 18241 46961 18269 46989
rect 18303 46961 18331 46989
rect 18117 38147 18145 38175
rect 18179 38147 18207 38175
rect 18241 38147 18269 38175
rect 18303 38147 18331 38175
rect 18117 38085 18145 38113
rect 18179 38085 18207 38113
rect 18241 38085 18269 38113
rect 18303 38085 18331 38113
rect 18117 38023 18145 38051
rect 18179 38023 18207 38051
rect 18241 38023 18269 38051
rect 18303 38023 18331 38051
rect 18117 37961 18145 37989
rect 18179 37961 18207 37989
rect 18241 37961 18269 37989
rect 18303 37961 18331 37989
rect 18117 29147 18145 29175
rect 18179 29147 18207 29175
rect 18241 29147 18269 29175
rect 18303 29147 18331 29175
rect 18117 29085 18145 29113
rect 18179 29085 18207 29113
rect 18241 29085 18269 29113
rect 18303 29085 18331 29113
rect 18117 29023 18145 29051
rect 18179 29023 18207 29051
rect 18241 29023 18269 29051
rect 18303 29023 18331 29051
rect 18117 28961 18145 28989
rect 18179 28961 18207 28989
rect 18241 28961 18269 28989
rect 18303 28961 18331 28989
rect 18117 20147 18145 20175
rect 18179 20147 18207 20175
rect 18241 20147 18269 20175
rect 18303 20147 18331 20175
rect 18117 20085 18145 20113
rect 18179 20085 18207 20113
rect 18241 20085 18269 20113
rect 18303 20085 18331 20113
rect 18117 20023 18145 20051
rect 18179 20023 18207 20051
rect 18241 20023 18269 20051
rect 18303 20023 18331 20051
rect 18117 19961 18145 19989
rect 18179 19961 18207 19989
rect 18241 19961 18269 19989
rect 18303 19961 18331 19989
rect 18117 11147 18145 11175
rect 18179 11147 18207 11175
rect 18241 11147 18269 11175
rect 18303 11147 18331 11175
rect 18117 11085 18145 11113
rect 18179 11085 18207 11113
rect 18241 11085 18269 11113
rect 18303 11085 18331 11113
rect 18117 11023 18145 11051
rect 18179 11023 18207 11051
rect 18241 11023 18269 11051
rect 18303 11023 18331 11051
rect 18117 10961 18145 10989
rect 18179 10961 18207 10989
rect 18241 10961 18269 10989
rect 18303 10961 18331 10989
rect 18117 2147 18145 2175
rect 18179 2147 18207 2175
rect 18241 2147 18269 2175
rect 18303 2147 18331 2175
rect 18117 2085 18145 2113
rect 18179 2085 18207 2113
rect 18241 2085 18269 2113
rect 18303 2085 18331 2113
rect 18117 2023 18145 2051
rect 18179 2023 18207 2051
rect 18241 2023 18269 2051
rect 18303 2023 18331 2051
rect 18117 1961 18145 1989
rect 18179 1961 18207 1989
rect 18241 1961 18269 1989
rect 18303 1961 18331 1989
rect 18117 -108 18145 -80
rect 18179 -108 18207 -80
rect 18241 -108 18269 -80
rect 18303 -108 18331 -80
rect 18117 -170 18145 -142
rect 18179 -170 18207 -142
rect 18241 -170 18269 -142
rect 18303 -170 18331 -142
rect 18117 -232 18145 -204
rect 18179 -232 18207 -204
rect 18241 -232 18269 -204
rect 18303 -232 18331 -204
rect 18117 -294 18145 -266
rect 18179 -294 18207 -266
rect 18241 -294 18269 -266
rect 18303 -294 18331 -266
rect 19977 299058 20005 299086
rect 20039 299058 20067 299086
rect 20101 299058 20129 299086
rect 20163 299058 20191 299086
rect 19977 298996 20005 299024
rect 20039 298996 20067 299024
rect 20101 298996 20129 299024
rect 20163 298996 20191 299024
rect 19977 298934 20005 298962
rect 20039 298934 20067 298962
rect 20101 298934 20129 298962
rect 20163 298934 20191 298962
rect 19977 298872 20005 298900
rect 20039 298872 20067 298900
rect 20101 298872 20129 298900
rect 20163 298872 20191 298900
rect 19977 293147 20005 293175
rect 20039 293147 20067 293175
rect 20101 293147 20129 293175
rect 20163 293147 20191 293175
rect 19977 293085 20005 293113
rect 20039 293085 20067 293113
rect 20101 293085 20129 293113
rect 20163 293085 20191 293113
rect 19977 293023 20005 293051
rect 20039 293023 20067 293051
rect 20101 293023 20129 293051
rect 20163 293023 20191 293051
rect 19977 292961 20005 292989
rect 20039 292961 20067 292989
rect 20101 292961 20129 292989
rect 20163 292961 20191 292989
rect 19977 284147 20005 284175
rect 20039 284147 20067 284175
rect 20101 284147 20129 284175
rect 20163 284147 20191 284175
rect 19977 284085 20005 284113
rect 20039 284085 20067 284113
rect 20101 284085 20129 284113
rect 20163 284085 20191 284113
rect 19977 284023 20005 284051
rect 20039 284023 20067 284051
rect 20101 284023 20129 284051
rect 20163 284023 20191 284051
rect 19977 283961 20005 283989
rect 20039 283961 20067 283989
rect 20101 283961 20129 283989
rect 20163 283961 20191 283989
rect 19977 275147 20005 275175
rect 20039 275147 20067 275175
rect 20101 275147 20129 275175
rect 20163 275147 20191 275175
rect 19977 275085 20005 275113
rect 20039 275085 20067 275113
rect 20101 275085 20129 275113
rect 20163 275085 20191 275113
rect 19977 275023 20005 275051
rect 20039 275023 20067 275051
rect 20101 275023 20129 275051
rect 20163 275023 20191 275051
rect 19977 274961 20005 274989
rect 20039 274961 20067 274989
rect 20101 274961 20129 274989
rect 20163 274961 20191 274989
rect 19977 266147 20005 266175
rect 20039 266147 20067 266175
rect 20101 266147 20129 266175
rect 20163 266147 20191 266175
rect 19977 266085 20005 266113
rect 20039 266085 20067 266113
rect 20101 266085 20129 266113
rect 20163 266085 20191 266113
rect 19977 266023 20005 266051
rect 20039 266023 20067 266051
rect 20101 266023 20129 266051
rect 20163 266023 20191 266051
rect 19977 265961 20005 265989
rect 20039 265961 20067 265989
rect 20101 265961 20129 265989
rect 20163 265961 20191 265989
rect 19977 257147 20005 257175
rect 20039 257147 20067 257175
rect 20101 257147 20129 257175
rect 20163 257147 20191 257175
rect 19977 257085 20005 257113
rect 20039 257085 20067 257113
rect 20101 257085 20129 257113
rect 20163 257085 20191 257113
rect 19977 257023 20005 257051
rect 20039 257023 20067 257051
rect 20101 257023 20129 257051
rect 20163 257023 20191 257051
rect 19977 256961 20005 256989
rect 20039 256961 20067 256989
rect 20101 256961 20129 256989
rect 20163 256961 20191 256989
rect 19977 248147 20005 248175
rect 20039 248147 20067 248175
rect 20101 248147 20129 248175
rect 20163 248147 20191 248175
rect 19977 248085 20005 248113
rect 20039 248085 20067 248113
rect 20101 248085 20129 248113
rect 20163 248085 20191 248113
rect 19977 248023 20005 248051
rect 20039 248023 20067 248051
rect 20101 248023 20129 248051
rect 20163 248023 20191 248051
rect 19977 247961 20005 247989
rect 20039 247961 20067 247989
rect 20101 247961 20129 247989
rect 20163 247961 20191 247989
rect 19977 239147 20005 239175
rect 20039 239147 20067 239175
rect 20101 239147 20129 239175
rect 20163 239147 20191 239175
rect 19977 239085 20005 239113
rect 20039 239085 20067 239113
rect 20101 239085 20129 239113
rect 20163 239085 20191 239113
rect 19977 239023 20005 239051
rect 20039 239023 20067 239051
rect 20101 239023 20129 239051
rect 20163 239023 20191 239051
rect 19977 238961 20005 238989
rect 20039 238961 20067 238989
rect 20101 238961 20129 238989
rect 20163 238961 20191 238989
rect 19977 230147 20005 230175
rect 20039 230147 20067 230175
rect 20101 230147 20129 230175
rect 20163 230147 20191 230175
rect 19977 230085 20005 230113
rect 20039 230085 20067 230113
rect 20101 230085 20129 230113
rect 20163 230085 20191 230113
rect 19977 230023 20005 230051
rect 20039 230023 20067 230051
rect 20101 230023 20129 230051
rect 20163 230023 20191 230051
rect 19977 229961 20005 229989
rect 20039 229961 20067 229989
rect 20101 229961 20129 229989
rect 20163 229961 20191 229989
rect 19977 221147 20005 221175
rect 20039 221147 20067 221175
rect 20101 221147 20129 221175
rect 20163 221147 20191 221175
rect 19977 221085 20005 221113
rect 20039 221085 20067 221113
rect 20101 221085 20129 221113
rect 20163 221085 20191 221113
rect 19977 221023 20005 221051
rect 20039 221023 20067 221051
rect 20101 221023 20129 221051
rect 20163 221023 20191 221051
rect 19977 220961 20005 220989
rect 20039 220961 20067 220989
rect 20101 220961 20129 220989
rect 20163 220961 20191 220989
rect 19977 212147 20005 212175
rect 20039 212147 20067 212175
rect 20101 212147 20129 212175
rect 20163 212147 20191 212175
rect 19977 212085 20005 212113
rect 20039 212085 20067 212113
rect 20101 212085 20129 212113
rect 20163 212085 20191 212113
rect 19977 212023 20005 212051
rect 20039 212023 20067 212051
rect 20101 212023 20129 212051
rect 20163 212023 20191 212051
rect 19977 211961 20005 211989
rect 20039 211961 20067 211989
rect 20101 211961 20129 211989
rect 20163 211961 20191 211989
rect 19977 203147 20005 203175
rect 20039 203147 20067 203175
rect 20101 203147 20129 203175
rect 20163 203147 20191 203175
rect 19977 203085 20005 203113
rect 20039 203085 20067 203113
rect 20101 203085 20129 203113
rect 20163 203085 20191 203113
rect 19977 203023 20005 203051
rect 20039 203023 20067 203051
rect 20101 203023 20129 203051
rect 20163 203023 20191 203051
rect 19977 202961 20005 202989
rect 20039 202961 20067 202989
rect 20101 202961 20129 202989
rect 20163 202961 20191 202989
rect 19977 194147 20005 194175
rect 20039 194147 20067 194175
rect 20101 194147 20129 194175
rect 20163 194147 20191 194175
rect 19977 194085 20005 194113
rect 20039 194085 20067 194113
rect 20101 194085 20129 194113
rect 20163 194085 20191 194113
rect 19977 194023 20005 194051
rect 20039 194023 20067 194051
rect 20101 194023 20129 194051
rect 20163 194023 20191 194051
rect 19977 193961 20005 193989
rect 20039 193961 20067 193989
rect 20101 193961 20129 193989
rect 20163 193961 20191 193989
rect 19977 185147 20005 185175
rect 20039 185147 20067 185175
rect 20101 185147 20129 185175
rect 20163 185147 20191 185175
rect 19977 185085 20005 185113
rect 20039 185085 20067 185113
rect 20101 185085 20129 185113
rect 20163 185085 20191 185113
rect 19977 185023 20005 185051
rect 20039 185023 20067 185051
rect 20101 185023 20129 185051
rect 20163 185023 20191 185051
rect 19977 184961 20005 184989
rect 20039 184961 20067 184989
rect 20101 184961 20129 184989
rect 20163 184961 20191 184989
rect 19977 176147 20005 176175
rect 20039 176147 20067 176175
rect 20101 176147 20129 176175
rect 20163 176147 20191 176175
rect 19977 176085 20005 176113
rect 20039 176085 20067 176113
rect 20101 176085 20129 176113
rect 20163 176085 20191 176113
rect 19977 176023 20005 176051
rect 20039 176023 20067 176051
rect 20101 176023 20129 176051
rect 20163 176023 20191 176051
rect 19977 175961 20005 175989
rect 20039 175961 20067 175989
rect 20101 175961 20129 175989
rect 20163 175961 20191 175989
rect 19977 167147 20005 167175
rect 20039 167147 20067 167175
rect 20101 167147 20129 167175
rect 20163 167147 20191 167175
rect 19977 167085 20005 167113
rect 20039 167085 20067 167113
rect 20101 167085 20129 167113
rect 20163 167085 20191 167113
rect 19977 167023 20005 167051
rect 20039 167023 20067 167051
rect 20101 167023 20129 167051
rect 20163 167023 20191 167051
rect 19977 166961 20005 166989
rect 20039 166961 20067 166989
rect 20101 166961 20129 166989
rect 20163 166961 20191 166989
rect 19977 158147 20005 158175
rect 20039 158147 20067 158175
rect 20101 158147 20129 158175
rect 20163 158147 20191 158175
rect 19977 158085 20005 158113
rect 20039 158085 20067 158113
rect 20101 158085 20129 158113
rect 20163 158085 20191 158113
rect 19977 158023 20005 158051
rect 20039 158023 20067 158051
rect 20101 158023 20129 158051
rect 20163 158023 20191 158051
rect 19977 157961 20005 157989
rect 20039 157961 20067 157989
rect 20101 157961 20129 157989
rect 20163 157961 20191 157989
rect 19977 149147 20005 149175
rect 20039 149147 20067 149175
rect 20101 149147 20129 149175
rect 20163 149147 20191 149175
rect 19977 149085 20005 149113
rect 20039 149085 20067 149113
rect 20101 149085 20129 149113
rect 20163 149085 20191 149113
rect 19977 149023 20005 149051
rect 20039 149023 20067 149051
rect 20101 149023 20129 149051
rect 20163 149023 20191 149051
rect 19977 148961 20005 148989
rect 20039 148961 20067 148989
rect 20101 148961 20129 148989
rect 20163 148961 20191 148989
rect 19977 140147 20005 140175
rect 20039 140147 20067 140175
rect 20101 140147 20129 140175
rect 20163 140147 20191 140175
rect 19977 140085 20005 140113
rect 20039 140085 20067 140113
rect 20101 140085 20129 140113
rect 20163 140085 20191 140113
rect 19977 140023 20005 140051
rect 20039 140023 20067 140051
rect 20101 140023 20129 140051
rect 20163 140023 20191 140051
rect 19977 139961 20005 139989
rect 20039 139961 20067 139989
rect 20101 139961 20129 139989
rect 20163 139961 20191 139989
rect 19977 131147 20005 131175
rect 20039 131147 20067 131175
rect 20101 131147 20129 131175
rect 20163 131147 20191 131175
rect 19977 131085 20005 131113
rect 20039 131085 20067 131113
rect 20101 131085 20129 131113
rect 20163 131085 20191 131113
rect 19977 131023 20005 131051
rect 20039 131023 20067 131051
rect 20101 131023 20129 131051
rect 20163 131023 20191 131051
rect 19977 130961 20005 130989
rect 20039 130961 20067 130989
rect 20101 130961 20129 130989
rect 20163 130961 20191 130989
rect 19977 122147 20005 122175
rect 20039 122147 20067 122175
rect 20101 122147 20129 122175
rect 20163 122147 20191 122175
rect 19977 122085 20005 122113
rect 20039 122085 20067 122113
rect 20101 122085 20129 122113
rect 20163 122085 20191 122113
rect 19977 122023 20005 122051
rect 20039 122023 20067 122051
rect 20101 122023 20129 122051
rect 20163 122023 20191 122051
rect 19977 121961 20005 121989
rect 20039 121961 20067 121989
rect 20101 121961 20129 121989
rect 20163 121961 20191 121989
rect 19977 113147 20005 113175
rect 20039 113147 20067 113175
rect 20101 113147 20129 113175
rect 20163 113147 20191 113175
rect 19977 113085 20005 113113
rect 20039 113085 20067 113113
rect 20101 113085 20129 113113
rect 20163 113085 20191 113113
rect 19977 113023 20005 113051
rect 20039 113023 20067 113051
rect 20101 113023 20129 113051
rect 20163 113023 20191 113051
rect 19977 112961 20005 112989
rect 20039 112961 20067 112989
rect 20101 112961 20129 112989
rect 20163 112961 20191 112989
rect 19977 104147 20005 104175
rect 20039 104147 20067 104175
rect 20101 104147 20129 104175
rect 20163 104147 20191 104175
rect 19977 104085 20005 104113
rect 20039 104085 20067 104113
rect 20101 104085 20129 104113
rect 20163 104085 20191 104113
rect 19977 104023 20005 104051
rect 20039 104023 20067 104051
rect 20101 104023 20129 104051
rect 20163 104023 20191 104051
rect 19977 103961 20005 103989
rect 20039 103961 20067 103989
rect 20101 103961 20129 103989
rect 20163 103961 20191 103989
rect 19977 95147 20005 95175
rect 20039 95147 20067 95175
rect 20101 95147 20129 95175
rect 20163 95147 20191 95175
rect 19977 95085 20005 95113
rect 20039 95085 20067 95113
rect 20101 95085 20129 95113
rect 20163 95085 20191 95113
rect 19977 95023 20005 95051
rect 20039 95023 20067 95051
rect 20101 95023 20129 95051
rect 20163 95023 20191 95051
rect 19977 94961 20005 94989
rect 20039 94961 20067 94989
rect 20101 94961 20129 94989
rect 20163 94961 20191 94989
rect 19977 86147 20005 86175
rect 20039 86147 20067 86175
rect 20101 86147 20129 86175
rect 20163 86147 20191 86175
rect 19977 86085 20005 86113
rect 20039 86085 20067 86113
rect 20101 86085 20129 86113
rect 20163 86085 20191 86113
rect 19977 86023 20005 86051
rect 20039 86023 20067 86051
rect 20101 86023 20129 86051
rect 20163 86023 20191 86051
rect 19977 85961 20005 85989
rect 20039 85961 20067 85989
rect 20101 85961 20129 85989
rect 20163 85961 20191 85989
rect 19977 77147 20005 77175
rect 20039 77147 20067 77175
rect 20101 77147 20129 77175
rect 20163 77147 20191 77175
rect 19977 77085 20005 77113
rect 20039 77085 20067 77113
rect 20101 77085 20129 77113
rect 20163 77085 20191 77113
rect 19977 77023 20005 77051
rect 20039 77023 20067 77051
rect 20101 77023 20129 77051
rect 20163 77023 20191 77051
rect 19977 76961 20005 76989
rect 20039 76961 20067 76989
rect 20101 76961 20129 76989
rect 20163 76961 20191 76989
rect 19977 68147 20005 68175
rect 20039 68147 20067 68175
rect 20101 68147 20129 68175
rect 20163 68147 20191 68175
rect 19977 68085 20005 68113
rect 20039 68085 20067 68113
rect 20101 68085 20129 68113
rect 20163 68085 20191 68113
rect 19977 68023 20005 68051
rect 20039 68023 20067 68051
rect 20101 68023 20129 68051
rect 20163 68023 20191 68051
rect 19977 67961 20005 67989
rect 20039 67961 20067 67989
rect 20101 67961 20129 67989
rect 20163 67961 20191 67989
rect 19977 59147 20005 59175
rect 20039 59147 20067 59175
rect 20101 59147 20129 59175
rect 20163 59147 20191 59175
rect 19977 59085 20005 59113
rect 20039 59085 20067 59113
rect 20101 59085 20129 59113
rect 20163 59085 20191 59113
rect 19977 59023 20005 59051
rect 20039 59023 20067 59051
rect 20101 59023 20129 59051
rect 20163 59023 20191 59051
rect 19977 58961 20005 58989
rect 20039 58961 20067 58989
rect 20101 58961 20129 58989
rect 20163 58961 20191 58989
rect 19977 50147 20005 50175
rect 20039 50147 20067 50175
rect 20101 50147 20129 50175
rect 20163 50147 20191 50175
rect 19977 50085 20005 50113
rect 20039 50085 20067 50113
rect 20101 50085 20129 50113
rect 20163 50085 20191 50113
rect 19977 50023 20005 50051
rect 20039 50023 20067 50051
rect 20101 50023 20129 50051
rect 20163 50023 20191 50051
rect 19977 49961 20005 49989
rect 20039 49961 20067 49989
rect 20101 49961 20129 49989
rect 20163 49961 20191 49989
rect 19977 41147 20005 41175
rect 20039 41147 20067 41175
rect 20101 41147 20129 41175
rect 20163 41147 20191 41175
rect 19977 41085 20005 41113
rect 20039 41085 20067 41113
rect 20101 41085 20129 41113
rect 20163 41085 20191 41113
rect 19977 41023 20005 41051
rect 20039 41023 20067 41051
rect 20101 41023 20129 41051
rect 20163 41023 20191 41051
rect 19977 40961 20005 40989
rect 20039 40961 20067 40989
rect 20101 40961 20129 40989
rect 20163 40961 20191 40989
rect 19977 32147 20005 32175
rect 20039 32147 20067 32175
rect 20101 32147 20129 32175
rect 20163 32147 20191 32175
rect 19977 32085 20005 32113
rect 20039 32085 20067 32113
rect 20101 32085 20129 32113
rect 20163 32085 20191 32113
rect 19977 32023 20005 32051
rect 20039 32023 20067 32051
rect 20101 32023 20129 32051
rect 20163 32023 20191 32051
rect 19977 31961 20005 31989
rect 20039 31961 20067 31989
rect 20101 31961 20129 31989
rect 20163 31961 20191 31989
rect 19977 23147 20005 23175
rect 20039 23147 20067 23175
rect 20101 23147 20129 23175
rect 20163 23147 20191 23175
rect 19977 23085 20005 23113
rect 20039 23085 20067 23113
rect 20101 23085 20129 23113
rect 20163 23085 20191 23113
rect 19977 23023 20005 23051
rect 20039 23023 20067 23051
rect 20101 23023 20129 23051
rect 20163 23023 20191 23051
rect 19977 22961 20005 22989
rect 20039 22961 20067 22989
rect 20101 22961 20129 22989
rect 20163 22961 20191 22989
rect 19977 14147 20005 14175
rect 20039 14147 20067 14175
rect 20101 14147 20129 14175
rect 20163 14147 20191 14175
rect 19977 14085 20005 14113
rect 20039 14085 20067 14113
rect 20101 14085 20129 14113
rect 20163 14085 20191 14113
rect 19977 14023 20005 14051
rect 20039 14023 20067 14051
rect 20101 14023 20129 14051
rect 20163 14023 20191 14051
rect 19977 13961 20005 13989
rect 20039 13961 20067 13989
rect 20101 13961 20129 13989
rect 20163 13961 20191 13989
rect 19977 5147 20005 5175
rect 20039 5147 20067 5175
rect 20101 5147 20129 5175
rect 20163 5147 20191 5175
rect 19977 5085 20005 5113
rect 20039 5085 20067 5113
rect 20101 5085 20129 5113
rect 20163 5085 20191 5113
rect 19977 5023 20005 5051
rect 20039 5023 20067 5051
rect 20101 5023 20129 5051
rect 20163 5023 20191 5051
rect 19977 4961 20005 4989
rect 20039 4961 20067 4989
rect 20101 4961 20129 4989
rect 20163 4961 20191 4989
rect 19977 -588 20005 -560
rect 20039 -588 20067 -560
rect 20101 -588 20129 -560
rect 20163 -588 20191 -560
rect 19977 -650 20005 -622
rect 20039 -650 20067 -622
rect 20101 -650 20129 -622
rect 20163 -650 20191 -622
rect 19977 -712 20005 -684
rect 20039 -712 20067 -684
rect 20101 -712 20129 -684
rect 20163 -712 20191 -684
rect 19977 -774 20005 -746
rect 20039 -774 20067 -746
rect 20101 -774 20129 -746
rect 20163 -774 20191 -746
rect 33477 298578 33505 298606
rect 33539 298578 33567 298606
rect 33601 298578 33629 298606
rect 33663 298578 33691 298606
rect 33477 298516 33505 298544
rect 33539 298516 33567 298544
rect 33601 298516 33629 298544
rect 33663 298516 33691 298544
rect 33477 298454 33505 298482
rect 33539 298454 33567 298482
rect 33601 298454 33629 298482
rect 33663 298454 33691 298482
rect 33477 298392 33505 298420
rect 33539 298392 33567 298420
rect 33601 298392 33629 298420
rect 33663 298392 33691 298420
rect 33477 290147 33505 290175
rect 33539 290147 33567 290175
rect 33601 290147 33629 290175
rect 33663 290147 33691 290175
rect 33477 290085 33505 290113
rect 33539 290085 33567 290113
rect 33601 290085 33629 290113
rect 33663 290085 33691 290113
rect 33477 290023 33505 290051
rect 33539 290023 33567 290051
rect 33601 290023 33629 290051
rect 33663 290023 33691 290051
rect 33477 289961 33505 289989
rect 33539 289961 33567 289989
rect 33601 289961 33629 289989
rect 33663 289961 33691 289989
rect 33477 281147 33505 281175
rect 33539 281147 33567 281175
rect 33601 281147 33629 281175
rect 33663 281147 33691 281175
rect 33477 281085 33505 281113
rect 33539 281085 33567 281113
rect 33601 281085 33629 281113
rect 33663 281085 33691 281113
rect 33477 281023 33505 281051
rect 33539 281023 33567 281051
rect 33601 281023 33629 281051
rect 33663 281023 33691 281051
rect 33477 280961 33505 280989
rect 33539 280961 33567 280989
rect 33601 280961 33629 280989
rect 33663 280961 33691 280989
rect 33477 272147 33505 272175
rect 33539 272147 33567 272175
rect 33601 272147 33629 272175
rect 33663 272147 33691 272175
rect 33477 272085 33505 272113
rect 33539 272085 33567 272113
rect 33601 272085 33629 272113
rect 33663 272085 33691 272113
rect 33477 272023 33505 272051
rect 33539 272023 33567 272051
rect 33601 272023 33629 272051
rect 33663 272023 33691 272051
rect 33477 271961 33505 271989
rect 33539 271961 33567 271989
rect 33601 271961 33629 271989
rect 33663 271961 33691 271989
rect 33477 263147 33505 263175
rect 33539 263147 33567 263175
rect 33601 263147 33629 263175
rect 33663 263147 33691 263175
rect 33477 263085 33505 263113
rect 33539 263085 33567 263113
rect 33601 263085 33629 263113
rect 33663 263085 33691 263113
rect 33477 263023 33505 263051
rect 33539 263023 33567 263051
rect 33601 263023 33629 263051
rect 33663 263023 33691 263051
rect 33477 262961 33505 262989
rect 33539 262961 33567 262989
rect 33601 262961 33629 262989
rect 33663 262961 33691 262989
rect 33477 254147 33505 254175
rect 33539 254147 33567 254175
rect 33601 254147 33629 254175
rect 33663 254147 33691 254175
rect 33477 254085 33505 254113
rect 33539 254085 33567 254113
rect 33601 254085 33629 254113
rect 33663 254085 33691 254113
rect 33477 254023 33505 254051
rect 33539 254023 33567 254051
rect 33601 254023 33629 254051
rect 33663 254023 33691 254051
rect 33477 253961 33505 253989
rect 33539 253961 33567 253989
rect 33601 253961 33629 253989
rect 33663 253961 33691 253989
rect 33477 245147 33505 245175
rect 33539 245147 33567 245175
rect 33601 245147 33629 245175
rect 33663 245147 33691 245175
rect 33477 245085 33505 245113
rect 33539 245085 33567 245113
rect 33601 245085 33629 245113
rect 33663 245085 33691 245113
rect 33477 245023 33505 245051
rect 33539 245023 33567 245051
rect 33601 245023 33629 245051
rect 33663 245023 33691 245051
rect 33477 244961 33505 244989
rect 33539 244961 33567 244989
rect 33601 244961 33629 244989
rect 33663 244961 33691 244989
rect 33477 236147 33505 236175
rect 33539 236147 33567 236175
rect 33601 236147 33629 236175
rect 33663 236147 33691 236175
rect 33477 236085 33505 236113
rect 33539 236085 33567 236113
rect 33601 236085 33629 236113
rect 33663 236085 33691 236113
rect 33477 236023 33505 236051
rect 33539 236023 33567 236051
rect 33601 236023 33629 236051
rect 33663 236023 33691 236051
rect 33477 235961 33505 235989
rect 33539 235961 33567 235989
rect 33601 235961 33629 235989
rect 33663 235961 33691 235989
rect 33477 227147 33505 227175
rect 33539 227147 33567 227175
rect 33601 227147 33629 227175
rect 33663 227147 33691 227175
rect 33477 227085 33505 227113
rect 33539 227085 33567 227113
rect 33601 227085 33629 227113
rect 33663 227085 33691 227113
rect 33477 227023 33505 227051
rect 33539 227023 33567 227051
rect 33601 227023 33629 227051
rect 33663 227023 33691 227051
rect 33477 226961 33505 226989
rect 33539 226961 33567 226989
rect 33601 226961 33629 226989
rect 33663 226961 33691 226989
rect 33477 218147 33505 218175
rect 33539 218147 33567 218175
rect 33601 218147 33629 218175
rect 33663 218147 33691 218175
rect 33477 218085 33505 218113
rect 33539 218085 33567 218113
rect 33601 218085 33629 218113
rect 33663 218085 33691 218113
rect 33477 218023 33505 218051
rect 33539 218023 33567 218051
rect 33601 218023 33629 218051
rect 33663 218023 33691 218051
rect 33477 217961 33505 217989
rect 33539 217961 33567 217989
rect 33601 217961 33629 217989
rect 33663 217961 33691 217989
rect 33477 209147 33505 209175
rect 33539 209147 33567 209175
rect 33601 209147 33629 209175
rect 33663 209147 33691 209175
rect 33477 209085 33505 209113
rect 33539 209085 33567 209113
rect 33601 209085 33629 209113
rect 33663 209085 33691 209113
rect 33477 209023 33505 209051
rect 33539 209023 33567 209051
rect 33601 209023 33629 209051
rect 33663 209023 33691 209051
rect 33477 208961 33505 208989
rect 33539 208961 33567 208989
rect 33601 208961 33629 208989
rect 33663 208961 33691 208989
rect 33477 200147 33505 200175
rect 33539 200147 33567 200175
rect 33601 200147 33629 200175
rect 33663 200147 33691 200175
rect 33477 200085 33505 200113
rect 33539 200085 33567 200113
rect 33601 200085 33629 200113
rect 33663 200085 33691 200113
rect 33477 200023 33505 200051
rect 33539 200023 33567 200051
rect 33601 200023 33629 200051
rect 33663 200023 33691 200051
rect 33477 199961 33505 199989
rect 33539 199961 33567 199989
rect 33601 199961 33629 199989
rect 33663 199961 33691 199989
rect 33477 191147 33505 191175
rect 33539 191147 33567 191175
rect 33601 191147 33629 191175
rect 33663 191147 33691 191175
rect 33477 191085 33505 191113
rect 33539 191085 33567 191113
rect 33601 191085 33629 191113
rect 33663 191085 33691 191113
rect 33477 191023 33505 191051
rect 33539 191023 33567 191051
rect 33601 191023 33629 191051
rect 33663 191023 33691 191051
rect 33477 190961 33505 190989
rect 33539 190961 33567 190989
rect 33601 190961 33629 190989
rect 33663 190961 33691 190989
rect 33477 182147 33505 182175
rect 33539 182147 33567 182175
rect 33601 182147 33629 182175
rect 33663 182147 33691 182175
rect 33477 182085 33505 182113
rect 33539 182085 33567 182113
rect 33601 182085 33629 182113
rect 33663 182085 33691 182113
rect 33477 182023 33505 182051
rect 33539 182023 33567 182051
rect 33601 182023 33629 182051
rect 33663 182023 33691 182051
rect 33477 181961 33505 181989
rect 33539 181961 33567 181989
rect 33601 181961 33629 181989
rect 33663 181961 33691 181989
rect 33477 173147 33505 173175
rect 33539 173147 33567 173175
rect 33601 173147 33629 173175
rect 33663 173147 33691 173175
rect 33477 173085 33505 173113
rect 33539 173085 33567 173113
rect 33601 173085 33629 173113
rect 33663 173085 33691 173113
rect 33477 173023 33505 173051
rect 33539 173023 33567 173051
rect 33601 173023 33629 173051
rect 33663 173023 33691 173051
rect 33477 172961 33505 172989
rect 33539 172961 33567 172989
rect 33601 172961 33629 172989
rect 33663 172961 33691 172989
rect 33477 164147 33505 164175
rect 33539 164147 33567 164175
rect 33601 164147 33629 164175
rect 33663 164147 33691 164175
rect 33477 164085 33505 164113
rect 33539 164085 33567 164113
rect 33601 164085 33629 164113
rect 33663 164085 33691 164113
rect 33477 164023 33505 164051
rect 33539 164023 33567 164051
rect 33601 164023 33629 164051
rect 33663 164023 33691 164051
rect 33477 163961 33505 163989
rect 33539 163961 33567 163989
rect 33601 163961 33629 163989
rect 33663 163961 33691 163989
rect 33477 155147 33505 155175
rect 33539 155147 33567 155175
rect 33601 155147 33629 155175
rect 33663 155147 33691 155175
rect 33477 155085 33505 155113
rect 33539 155085 33567 155113
rect 33601 155085 33629 155113
rect 33663 155085 33691 155113
rect 33477 155023 33505 155051
rect 33539 155023 33567 155051
rect 33601 155023 33629 155051
rect 33663 155023 33691 155051
rect 33477 154961 33505 154989
rect 33539 154961 33567 154989
rect 33601 154961 33629 154989
rect 33663 154961 33691 154989
rect 33477 146147 33505 146175
rect 33539 146147 33567 146175
rect 33601 146147 33629 146175
rect 33663 146147 33691 146175
rect 33477 146085 33505 146113
rect 33539 146085 33567 146113
rect 33601 146085 33629 146113
rect 33663 146085 33691 146113
rect 33477 146023 33505 146051
rect 33539 146023 33567 146051
rect 33601 146023 33629 146051
rect 33663 146023 33691 146051
rect 33477 145961 33505 145989
rect 33539 145961 33567 145989
rect 33601 145961 33629 145989
rect 33663 145961 33691 145989
rect 33477 137147 33505 137175
rect 33539 137147 33567 137175
rect 33601 137147 33629 137175
rect 33663 137147 33691 137175
rect 33477 137085 33505 137113
rect 33539 137085 33567 137113
rect 33601 137085 33629 137113
rect 33663 137085 33691 137113
rect 33477 137023 33505 137051
rect 33539 137023 33567 137051
rect 33601 137023 33629 137051
rect 33663 137023 33691 137051
rect 33477 136961 33505 136989
rect 33539 136961 33567 136989
rect 33601 136961 33629 136989
rect 33663 136961 33691 136989
rect 33477 128147 33505 128175
rect 33539 128147 33567 128175
rect 33601 128147 33629 128175
rect 33663 128147 33691 128175
rect 33477 128085 33505 128113
rect 33539 128085 33567 128113
rect 33601 128085 33629 128113
rect 33663 128085 33691 128113
rect 33477 128023 33505 128051
rect 33539 128023 33567 128051
rect 33601 128023 33629 128051
rect 33663 128023 33691 128051
rect 33477 127961 33505 127989
rect 33539 127961 33567 127989
rect 33601 127961 33629 127989
rect 33663 127961 33691 127989
rect 33477 119147 33505 119175
rect 33539 119147 33567 119175
rect 33601 119147 33629 119175
rect 33663 119147 33691 119175
rect 33477 119085 33505 119113
rect 33539 119085 33567 119113
rect 33601 119085 33629 119113
rect 33663 119085 33691 119113
rect 33477 119023 33505 119051
rect 33539 119023 33567 119051
rect 33601 119023 33629 119051
rect 33663 119023 33691 119051
rect 33477 118961 33505 118989
rect 33539 118961 33567 118989
rect 33601 118961 33629 118989
rect 33663 118961 33691 118989
rect 33477 110147 33505 110175
rect 33539 110147 33567 110175
rect 33601 110147 33629 110175
rect 33663 110147 33691 110175
rect 33477 110085 33505 110113
rect 33539 110085 33567 110113
rect 33601 110085 33629 110113
rect 33663 110085 33691 110113
rect 33477 110023 33505 110051
rect 33539 110023 33567 110051
rect 33601 110023 33629 110051
rect 33663 110023 33691 110051
rect 33477 109961 33505 109989
rect 33539 109961 33567 109989
rect 33601 109961 33629 109989
rect 33663 109961 33691 109989
rect 33477 101147 33505 101175
rect 33539 101147 33567 101175
rect 33601 101147 33629 101175
rect 33663 101147 33691 101175
rect 33477 101085 33505 101113
rect 33539 101085 33567 101113
rect 33601 101085 33629 101113
rect 33663 101085 33691 101113
rect 33477 101023 33505 101051
rect 33539 101023 33567 101051
rect 33601 101023 33629 101051
rect 33663 101023 33691 101051
rect 33477 100961 33505 100989
rect 33539 100961 33567 100989
rect 33601 100961 33629 100989
rect 33663 100961 33691 100989
rect 33477 92147 33505 92175
rect 33539 92147 33567 92175
rect 33601 92147 33629 92175
rect 33663 92147 33691 92175
rect 33477 92085 33505 92113
rect 33539 92085 33567 92113
rect 33601 92085 33629 92113
rect 33663 92085 33691 92113
rect 33477 92023 33505 92051
rect 33539 92023 33567 92051
rect 33601 92023 33629 92051
rect 33663 92023 33691 92051
rect 33477 91961 33505 91989
rect 33539 91961 33567 91989
rect 33601 91961 33629 91989
rect 33663 91961 33691 91989
rect 33477 83147 33505 83175
rect 33539 83147 33567 83175
rect 33601 83147 33629 83175
rect 33663 83147 33691 83175
rect 33477 83085 33505 83113
rect 33539 83085 33567 83113
rect 33601 83085 33629 83113
rect 33663 83085 33691 83113
rect 33477 83023 33505 83051
rect 33539 83023 33567 83051
rect 33601 83023 33629 83051
rect 33663 83023 33691 83051
rect 33477 82961 33505 82989
rect 33539 82961 33567 82989
rect 33601 82961 33629 82989
rect 33663 82961 33691 82989
rect 33477 74147 33505 74175
rect 33539 74147 33567 74175
rect 33601 74147 33629 74175
rect 33663 74147 33691 74175
rect 33477 74085 33505 74113
rect 33539 74085 33567 74113
rect 33601 74085 33629 74113
rect 33663 74085 33691 74113
rect 33477 74023 33505 74051
rect 33539 74023 33567 74051
rect 33601 74023 33629 74051
rect 33663 74023 33691 74051
rect 33477 73961 33505 73989
rect 33539 73961 33567 73989
rect 33601 73961 33629 73989
rect 33663 73961 33691 73989
rect 33477 65147 33505 65175
rect 33539 65147 33567 65175
rect 33601 65147 33629 65175
rect 33663 65147 33691 65175
rect 33477 65085 33505 65113
rect 33539 65085 33567 65113
rect 33601 65085 33629 65113
rect 33663 65085 33691 65113
rect 33477 65023 33505 65051
rect 33539 65023 33567 65051
rect 33601 65023 33629 65051
rect 33663 65023 33691 65051
rect 33477 64961 33505 64989
rect 33539 64961 33567 64989
rect 33601 64961 33629 64989
rect 33663 64961 33691 64989
rect 33477 56147 33505 56175
rect 33539 56147 33567 56175
rect 33601 56147 33629 56175
rect 33663 56147 33691 56175
rect 33477 56085 33505 56113
rect 33539 56085 33567 56113
rect 33601 56085 33629 56113
rect 33663 56085 33691 56113
rect 33477 56023 33505 56051
rect 33539 56023 33567 56051
rect 33601 56023 33629 56051
rect 33663 56023 33691 56051
rect 33477 55961 33505 55989
rect 33539 55961 33567 55989
rect 33601 55961 33629 55989
rect 33663 55961 33691 55989
rect 33477 47147 33505 47175
rect 33539 47147 33567 47175
rect 33601 47147 33629 47175
rect 33663 47147 33691 47175
rect 33477 47085 33505 47113
rect 33539 47085 33567 47113
rect 33601 47085 33629 47113
rect 33663 47085 33691 47113
rect 33477 47023 33505 47051
rect 33539 47023 33567 47051
rect 33601 47023 33629 47051
rect 33663 47023 33691 47051
rect 33477 46961 33505 46989
rect 33539 46961 33567 46989
rect 33601 46961 33629 46989
rect 33663 46961 33691 46989
rect 33477 38147 33505 38175
rect 33539 38147 33567 38175
rect 33601 38147 33629 38175
rect 33663 38147 33691 38175
rect 33477 38085 33505 38113
rect 33539 38085 33567 38113
rect 33601 38085 33629 38113
rect 33663 38085 33691 38113
rect 33477 38023 33505 38051
rect 33539 38023 33567 38051
rect 33601 38023 33629 38051
rect 33663 38023 33691 38051
rect 33477 37961 33505 37989
rect 33539 37961 33567 37989
rect 33601 37961 33629 37989
rect 33663 37961 33691 37989
rect 33477 29147 33505 29175
rect 33539 29147 33567 29175
rect 33601 29147 33629 29175
rect 33663 29147 33691 29175
rect 33477 29085 33505 29113
rect 33539 29085 33567 29113
rect 33601 29085 33629 29113
rect 33663 29085 33691 29113
rect 33477 29023 33505 29051
rect 33539 29023 33567 29051
rect 33601 29023 33629 29051
rect 33663 29023 33691 29051
rect 33477 28961 33505 28989
rect 33539 28961 33567 28989
rect 33601 28961 33629 28989
rect 33663 28961 33691 28989
rect 33477 20147 33505 20175
rect 33539 20147 33567 20175
rect 33601 20147 33629 20175
rect 33663 20147 33691 20175
rect 33477 20085 33505 20113
rect 33539 20085 33567 20113
rect 33601 20085 33629 20113
rect 33663 20085 33691 20113
rect 33477 20023 33505 20051
rect 33539 20023 33567 20051
rect 33601 20023 33629 20051
rect 33663 20023 33691 20051
rect 33477 19961 33505 19989
rect 33539 19961 33567 19989
rect 33601 19961 33629 19989
rect 33663 19961 33691 19989
rect 33477 11147 33505 11175
rect 33539 11147 33567 11175
rect 33601 11147 33629 11175
rect 33663 11147 33691 11175
rect 33477 11085 33505 11113
rect 33539 11085 33567 11113
rect 33601 11085 33629 11113
rect 33663 11085 33691 11113
rect 33477 11023 33505 11051
rect 33539 11023 33567 11051
rect 33601 11023 33629 11051
rect 33663 11023 33691 11051
rect 33477 10961 33505 10989
rect 33539 10961 33567 10989
rect 33601 10961 33629 10989
rect 33663 10961 33691 10989
rect 33477 2147 33505 2175
rect 33539 2147 33567 2175
rect 33601 2147 33629 2175
rect 33663 2147 33691 2175
rect 33477 2085 33505 2113
rect 33539 2085 33567 2113
rect 33601 2085 33629 2113
rect 33663 2085 33691 2113
rect 33477 2023 33505 2051
rect 33539 2023 33567 2051
rect 33601 2023 33629 2051
rect 33663 2023 33691 2051
rect 33477 1961 33505 1989
rect 33539 1961 33567 1989
rect 33601 1961 33629 1989
rect 33663 1961 33691 1989
rect 33477 -108 33505 -80
rect 33539 -108 33567 -80
rect 33601 -108 33629 -80
rect 33663 -108 33691 -80
rect 33477 -170 33505 -142
rect 33539 -170 33567 -142
rect 33601 -170 33629 -142
rect 33663 -170 33691 -142
rect 33477 -232 33505 -204
rect 33539 -232 33567 -204
rect 33601 -232 33629 -204
rect 33663 -232 33691 -204
rect 33477 -294 33505 -266
rect 33539 -294 33567 -266
rect 33601 -294 33629 -266
rect 33663 -294 33691 -266
rect 35337 299058 35365 299086
rect 35399 299058 35427 299086
rect 35461 299058 35489 299086
rect 35523 299058 35551 299086
rect 35337 298996 35365 299024
rect 35399 298996 35427 299024
rect 35461 298996 35489 299024
rect 35523 298996 35551 299024
rect 35337 298934 35365 298962
rect 35399 298934 35427 298962
rect 35461 298934 35489 298962
rect 35523 298934 35551 298962
rect 35337 298872 35365 298900
rect 35399 298872 35427 298900
rect 35461 298872 35489 298900
rect 35523 298872 35551 298900
rect 35337 293147 35365 293175
rect 35399 293147 35427 293175
rect 35461 293147 35489 293175
rect 35523 293147 35551 293175
rect 35337 293085 35365 293113
rect 35399 293085 35427 293113
rect 35461 293085 35489 293113
rect 35523 293085 35551 293113
rect 35337 293023 35365 293051
rect 35399 293023 35427 293051
rect 35461 293023 35489 293051
rect 35523 293023 35551 293051
rect 35337 292961 35365 292989
rect 35399 292961 35427 292989
rect 35461 292961 35489 292989
rect 35523 292961 35551 292989
rect 35337 284147 35365 284175
rect 35399 284147 35427 284175
rect 35461 284147 35489 284175
rect 35523 284147 35551 284175
rect 35337 284085 35365 284113
rect 35399 284085 35427 284113
rect 35461 284085 35489 284113
rect 35523 284085 35551 284113
rect 35337 284023 35365 284051
rect 35399 284023 35427 284051
rect 35461 284023 35489 284051
rect 35523 284023 35551 284051
rect 35337 283961 35365 283989
rect 35399 283961 35427 283989
rect 35461 283961 35489 283989
rect 35523 283961 35551 283989
rect 35337 275147 35365 275175
rect 35399 275147 35427 275175
rect 35461 275147 35489 275175
rect 35523 275147 35551 275175
rect 35337 275085 35365 275113
rect 35399 275085 35427 275113
rect 35461 275085 35489 275113
rect 35523 275085 35551 275113
rect 35337 275023 35365 275051
rect 35399 275023 35427 275051
rect 35461 275023 35489 275051
rect 35523 275023 35551 275051
rect 35337 274961 35365 274989
rect 35399 274961 35427 274989
rect 35461 274961 35489 274989
rect 35523 274961 35551 274989
rect 35337 266147 35365 266175
rect 35399 266147 35427 266175
rect 35461 266147 35489 266175
rect 35523 266147 35551 266175
rect 35337 266085 35365 266113
rect 35399 266085 35427 266113
rect 35461 266085 35489 266113
rect 35523 266085 35551 266113
rect 35337 266023 35365 266051
rect 35399 266023 35427 266051
rect 35461 266023 35489 266051
rect 35523 266023 35551 266051
rect 35337 265961 35365 265989
rect 35399 265961 35427 265989
rect 35461 265961 35489 265989
rect 35523 265961 35551 265989
rect 35337 257147 35365 257175
rect 35399 257147 35427 257175
rect 35461 257147 35489 257175
rect 35523 257147 35551 257175
rect 35337 257085 35365 257113
rect 35399 257085 35427 257113
rect 35461 257085 35489 257113
rect 35523 257085 35551 257113
rect 35337 257023 35365 257051
rect 35399 257023 35427 257051
rect 35461 257023 35489 257051
rect 35523 257023 35551 257051
rect 35337 256961 35365 256989
rect 35399 256961 35427 256989
rect 35461 256961 35489 256989
rect 35523 256961 35551 256989
rect 35337 248147 35365 248175
rect 35399 248147 35427 248175
rect 35461 248147 35489 248175
rect 35523 248147 35551 248175
rect 35337 248085 35365 248113
rect 35399 248085 35427 248113
rect 35461 248085 35489 248113
rect 35523 248085 35551 248113
rect 35337 248023 35365 248051
rect 35399 248023 35427 248051
rect 35461 248023 35489 248051
rect 35523 248023 35551 248051
rect 35337 247961 35365 247989
rect 35399 247961 35427 247989
rect 35461 247961 35489 247989
rect 35523 247961 35551 247989
rect 35337 239147 35365 239175
rect 35399 239147 35427 239175
rect 35461 239147 35489 239175
rect 35523 239147 35551 239175
rect 35337 239085 35365 239113
rect 35399 239085 35427 239113
rect 35461 239085 35489 239113
rect 35523 239085 35551 239113
rect 35337 239023 35365 239051
rect 35399 239023 35427 239051
rect 35461 239023 35489 239051
rect 35523 239023 35551 239051
rect 35337 238961 35365 238989
rect 35399 238961 35427 238989
rect 35461 238961 35489 238989
rect 35523 238961 35551 238989
rect 35337 230147 35365 230175
rect 35399 230147 35427 230175
rect 35461 230147 35489 230175
rect 35523 230147 35551 230175
rect 35337 230085 35365 230113
rect 35399 230085 35427 230113
rect 35461 230085 35489 230113
rect 35523 230085 35551 230113
rect 35337 230023 35365 230051
rect 35399 230023 35427 230051
rect 35461 230023 35489 230051
rect 35523 230023 35551 230051
rect 35337 229961 35365 229989
rect 35399 229961 35427 229989
rect 35461 229961 35489 229989
rect 35523 229961 35551 229989
rect 35337 221147 35365 221175
rect 35399 221147 35427 221175
rect 35461 221147 35489 221175
rect 35523 221147 35551 221175
rect 35337 221085 35365 221113
rect 35399 221085 35427 221113
rect 35461 221085 35489 221113
rect 35523 221085 35551 221113
rect 35337 221023 35365 221051
rect 35399 221023 35427 221051
rect 35461 221023 35489 221051
rect 35523 221023 35551 221051
rect 35337 220961 35365 220989
rect 35399 220961 35427 220989
rect 35461 220961 35489 220989
rect 35523 220961 35551 220989
rect 35337 212147 35365 212175
rect 35399 212147 35427 212175
rect 35461 212147 35489 212175
rect 35523 212147 35551 212175
rect 35337 212085 35365 212113
rect 35399 212085 35427 212113
rect 35461 212085 35489 212113
rect 35523 212085 35551 212113
rect 35337 212023 35365 212051
rect 35399 212023 35427 212051
rect 35461 212023 35489 212051
rect 35523 212023 35551 212051
rect 35337 211961 35365 211989
rect 35399 211961 35427 211989
rect 35461 211961 35489 211989
rect 35523 211961 35551 211989
rect 35337 203147 35365 203175
rect 35399 203147 35427 203175
rect 35461 203147 35489 203175
rect 35523 203147 35551 203175
rect 35337 203085 35365 203113
rect 35399 203085 35427 203113
rect 35461 203085 35489 203113
rect 35523 203085 35551 203113
rect 35337 203023 35365 203051
rect 35399 203023 35427 203051
rect 35461 203023 35489 203051
rect 35523 203023 35551 203051
rect 35337 202961 35365 202989
rect 35399 202961 35427 202989
rect 35461 202961 35489 202989
rect 35523 202961 35551 202989
rect 35337 194147 35365 194175
rect 35399 194147 35427 194175
rect 35461 194147 35489 194175
rect 35523 194147 35551 194175
rect 35337 194085 35365 194113
rect 35399 194085 35427 194113
rect 35461 194085 35489 194113
rect 35523 194085 35551 194113
rect 35337 194023 35365 194051
rect 35399 194023 35427 194051
rect 35461 194023 35489 194051
rect 35523 194023 35551 194051
rect 35337 193961 35365 193989
rect 35399 193961 35427 193989
rect 35461 193961 35489 193989
rect 35523 193961 35551 193989
rect 35337 185147 35365 185175
rect 35399 185147 35427 185175
rect 35461 185147 35489 185175
rect 35523 185147 35551 185175
rect 35337 185085 35365 185113
rect 35399 185085 35427 185113
rect 35461 185085 35489 185113
rect 35523 185085 35551 185113
rect 35337 185023 35365 185051
rect 35399 185023 35427 185051
rect 35461 185023 35489 185051
rect 35523 185023 35551 185051
rect 35337 184961 35365 184989
rect 35399 184961 35427 184989
rect 35461 184961 35489 184989
rect 35523 184961 35551 184989
rect 35337 176147 35365 176175
rect 35399 176147 35427 176175
rect 35461 176147 35489 176175
rect 35523 176147 35551 176175
rect 35337 176085 35365 176113
rect 35399 176085 35427 176113
rect 35461 176085 35489 176113
rect 35523 176085 35551 176113
rect 35337 176023 35365 176051
rect 35399 176023 35427 176051
rect 35461 176023 35489 176051
rect 35523 176023 35551 176051
rect 35337 175961 35365 175989
rect 35399 175961 35427 175989
rect 35461 175961 35489 175989
rect 35523 175961 35551 175989
rect 35337 167147 35365 167175
rect 35399 167147 35427 167175
rect 35461 167147 35489 167175
rect 35523 167147 35551 167175
rect 35337 167085 35365 167113
rect 35399 167085 35427 167113
rect 35461 167085 35489 167113
rect 35523 167085 35551 167113
rect 35337 167023 35365 167051
rect 35399 167023 35427 167051
rect 35461 167023 35489 167051
rect 35523 167023 35551 167051
rect 35337 166961 35365 166989
rect 35399 166961 35427 166989
rect 35461 166961 35489 166989
rect 35523 166961 35551 166989
rect 35337 158147 35365 158175
rect 35399 158147 35427 158175
rect 35461 158147 35489 158175
rect 35523 158147 35551 158175
rect 35337 158085 35365 158113
rect 35399 158085 35427 158113
rect 35461 158085 35489 158113
rect 35523 158085 35551 158113
rect 35337 158023 35365 158051
rect 35399 158023 35427 158051
rect 35461 158023 35489 158051
rect 35523 158023 35551 158051
rect 35337 157961 35365 157989
rect 35399 157961 35427 157989
rect 35461 157961 35489 157989
rect 35523 157961 35551 157989
rect 35337 149147 35365 149175
rect 35399 149147 35427 149175
rect 35461 149147 35489 149175
rect 35523 149147 35551 149175
rect 35337 149085 35365 149113
rect 35399 149085 35427 149113
rect 35461 149085 35489 149113
rect 35523 149085 35551 149113
rect 35337 149023 35365 149051
rect 35399 149023 35427 149051
rect 35461 149023 35489 149051
rect 35523 149023 35551 149051
rect 35337 148961 35365 148989
rect 35399 148961 35427 148989
rect 35461 148961 35489 148989
rect 35523 148961 35551 148989
rect 35337 140147 35365 140175
rect 35399 140147 35427 140175
rect 35461 140147 35489 140175
rect 35523 140147 35551 140175
rect 35337 140085 35365 140113
rect 35399 140085 35427 140113
rect 35461 140085 35489 140113
rect 35523 140085 35551 140113
rect 35337 140023 35365 140051
rect 35399 140023 35427 140051
rect 35461 140023 35489 140051
rect 35523 140023 35551 140051
rect 35337 139961 35365 139989
rect 35399 139961 35427 139989
rect 35461 139961 35489 139989
rect 35523 139961 35551 139989
rect 35337 131147 35365 131175
rect 35399 131147 35427 131175
rect 35461 131147 35489 131175
rect 35523 131147 35551 131175
rect 35337 131085 35365 131113
rect 35399 131085 35427 131113
rect 35461 131085 35489 131113
rect 35523 131085 35551 131113
rect 35337 131023 35365 131051
rect 35399 131023 35427 131051
rect 35461 131023 35489 131051
rect 35523 131023 35551 131051
rect 35337 130961 35365 130989
rect 35399 130961 35427 130989
rect 35461 130961 35489 130989
rect 35523 130961 35551 130989
rect 35337 122147 35365 122175
rect 35399 122147 35427 122175
rect 35461 122147 35489 122175
rect 35523 122147 35551 122175
rect 35337 122085 35365 122113
rect 35399 122085 35427 122113
rect 35461 122085 35489 122113
rect 35523 122085 35551 122113
rect 35337 122023 35365 122051
rect 35399 122023 35427 122051
rect 35461 122023 35489 122051
rect 35523 122023 35551 122051
rect 35337 121961 35365 121989
rect 35399 121961 35427 121989
rect 35461 121961 35489 121989
rect 35523 121961 35551 121989
rect 35337 113147 35365 113175
rect 35399 113147 35427 113175
rect 35461 113147 35489 113175
rect 35523 113147 35551 113175
rect 35337 113085 35365 113113
rect 35399 113085 35427 113113
rect 35461 113085 35489 113113
rect 35523 113085 35551 113113
rect 35337 113023 35365 113051
rect 35399 113023 35427 113051
rect 35461 113023 35489 113051
rect 35523 113023 35551 113051
rect 35337 112961 35365 112989
rect 35399 112961 35427 112989
rect 35461 112961 35489 112989
rect 35523 112961 35551 112989
rect 35337 104147 35365 104175
rect 35399 104147 35427 104175
rect 35461 104147 35489 104175
rect 35523 104147 35551 104175
rect 35337 104085 35365 104113
rect 35399 104085 35427 104113
rect 35461 104085 35489 104113
rect 35523 104085 35551 104113
rect 35337 104023 35365 104051
rect 35399 104023 35427 104051
rect 35461 104023 35489 104051
rect 35523 104023 35551 104051
rect 35337 103961 35365 103989
rect 35399 103961 35427 103989
rect 35461 103961 35489 103989
rect 35523 103961 35551 103989
rect 35337 95147 35365 95175
rect 35399 95147 35427 95175
rect 35461 95147 35489 95175
rect 35523 95147 35551 95175
rect 35337 95085 35365 95113
rect 35399 95085 35427 95113
rect 35461 95085 35489 95113
rect 35523 95085 35551 95113
rect 35337 95023 35365 95051
rect 35399 95023 35427 95051
rect 35461 95023 35489 95051
rect 35523 95023 35551 95051
rect 35337 94961 35365 94989
rect 35399 94961 35427 94989
rect 35461 94961 35489 94989
rect 35523 94961 35551 94989
rect 35337 86147 35365 86175
rect 35399 86147 35427 86175
rect 35461 86147 35489 86175
rect 35523 86147 35551 86175
rect 35337 86085 35365 86113
rect 35399 86085 35427 86113
rect 35461 86085 35489 86113
rect 35523 86085 35551 86113
rect 35337 86023 35365 86051
rect 35399 86023 35427 86051
rect 35461 86023 35489 86051
rect 35523 86023 35551 86051
rect 35337 85961 35365 85989
rect 35399 85961 35427 85989
rect 35461 85961 35489 85989
rect 35523 85961 35551 85989
rect 35337 77147 35365 77175
rect 35399 77147 35427 77175
rect 35461 77147 35489 77175
rect 35523 77147 35551 77175
rect 35337 77085 35365 77113
rect 35399 77085 35427 77113
rect 35461 77085 35489 77113
rect 35523 77085 35551 77113
rect 35337 77023 35365 77051
rect 35399 77023 35427 77051
rect 35461 77023 35489 77051
rect 35523 77023 35551 77051
rect 35337 76961 35365 76989
rect 35399 76961 35427 76989
rect 35461 76961 35489 76989
rect 35523 76961 35551 76989
rect 35337 68147 35365 68175
rect 35399 68147 35427 68175
rect 35461 68147 35489 68175
rect 35523 68147 35551 68175
rect 35337 68085 35365 68113
rect 35399 68085 35427 68113
rect 35461 68085 35489 68113
rect 35523 68085 35551 68113
rect 35337 68023 35365 68051
rect 35399 68023 35427 68051
rect 35461 68023 35489 68051
rect 35523 68023 35551 68051
rect 35337 67961 35365 67989
rect 35399 67961 35427 67989
rect 35461 67961 35489 67989
rect 35523 67961 35551 67989
rect 35337 59147 35365 59175
rect 35399 59147 35427 59175
rect 35461 59147 35489 59175
rect 35523 59147 35551 59175
rect 35337 59085 35365 59113
rect 35399 59085 35427 59113
rect 35461 59085 35489 59113
rect 35523 59085 35551 59113
rect 35337 59023 35365 59051
rect 35399 59023 35427 59051
rect 35461 59023 35489 59051
rect 35523 59023 35551 59051
rect 35337 58961 35365 58989
rect 35399 58961 35427 58989
rect 35461 58961 35489 58989
rect 35523 58961 35551 58989
rect 35337 50147 35365 50175
rect 35399 50147 35427 50175
rect 35461 50147 35489 50175
rect 35523 50147 35551 50175
rect 35337 50085 35365 50113
rect 35399 50085 35427 50113
rect 35461 50085 35489 50113
rect 35523 50085 35551 50113
rect 35337 50023 35365 50051
rect 35399 50023 35427 50051
rect 35461 50023 35489 50051
rect 35523 50023 35551 50051
rect 35337 49961 35365 49989
rect 35399 49961 35427 49989
rect 35461 49961 35489 49989
rect 35523 49961 35551 49989
rect 35337 41147 35365 41175
rect 35399 41147 35427 41175
rect 35461 41147 35489 41175
rect 35523 41147 35551 41175
rect 35337 41085 35365 41113
rect 35399 41085 35427 41113
rect 35461 41085 35489 41113
rect 35523 41085 35551 41113
rect 35337 41023 35365 41051
rect 35399 41023 35427 41051
rect 35461 41023 35489 41051
rect 35523 41023 35551 41051
rect 35337 40961 35365 40989
rect 35399 40961 35427 40989
rect 35461 40961 35489 40989
rect 35523 40961 35551 40989
rect 35337 32147 35365 32175
rect 35399 32147 35427 32175
rect 35461 32147 35489 32175
rect 35523 32147 35551 32175
rect 35337 32085 35365 32113
rect 35399 32085 35427 32113
rect 35461 32085 35489 32113
rect 35523 32085 35551 32113
rect 35337 32023 35365 32051
rect 35399 32023 35427 32051
rect 35461 32023 35489 32051
rect 35523 32023 35551 32051
rect 35337 31961 35365 31989
rect 35399 31961 35427 31989
rect 35461 31961 35489 31989
rect 35523 31961 35551 31989
rect 35337 23147 35365 23175
rect 35399 23147 35427 23175
rect 35461 23147 35489 23175
rect 35523 23147 35551 23175
rect 35337 23085 35365 23113
rect 35399 23085 35427 23113
rect 35461 23085 35489 23113
rect 35523 23085 35551 23113
rect 35337 23023 35365 23051
rect 35399 23023 35427 23051
rect 35461 23023 35489 23051
rect 35523 23023 35551 23051
rect 35337 22961 35365 22989
rect 35399 22961 35427 22989
rect 35461 22961 35489 22989
rect 35523 22961 35551 22989
rect 35337 14147 35365 14175
rect 35399 14147 35427 14175
rect 35461 14147 35489 14175
rect 35523 14147 35551 14175
rect 35337 14085 35365 14113
rect 35399 14085 35427 14113
rect 35461 14085 35489 14113
rect 35523 14085 35551 14113
rect 35337 14023 35365 14051
rect 35399 14023 35427 14051
rect 35461 14023 35489 14051
rect 35523 14023 35551 14051
rect 35337 13961 35365 13989
rect 35399 13961 35427 13989
rect 35461 13961 35489 13989
rect 35523 13961 35551 13989
rect 35337 5147 35365 5175
rect 35399 5147 35427 5175
rect 35461 5147 35489 5175
rect 35523 5147 35551 5175
rect 35337 5085 35365 5113
rect 35399 5085 35427 5113
rect 35461 5085 35489 5113
rect 35523 5085 35551 5113
rect 35337 5023 35365 5051
rect 35399 5023 35427 5051
rect 35461 5023 35489 5051
rect 35523 5023 35551 5051
rect 35337 4961 35365 4989
rect 35399 4961 35427 4989
rect 35461 4961 35489 4989
rect 35523 4961 35551 4989
rect 35337 -588 35365 -560
rect 35399 -588 35427 -560
rect 35461 -588 35489 -560
rect 35523 -588 35551 -560
rect 35337 -650 35365 -622
rect 35399 -650 35427 -622
rect 35461 -650 35489 -622
rect 35523 -650 35551 -622
rect 35337 -712 35365 -684
rect 35399 -712 35427 -684
rect 35461 -712 35489 -684
rect 35523 -712 35551 -684
rect 35337 -774 35365 -746
rect 35399 -774 35427 -746
rect 35461 -774 35489 -746
rect 35523 -774 35551 -746
rect 48837 298578 48865 298606
rect 48899 298578 48927 298606
rect 48961 298578 48989 298606
rect 49023 298578 49051 298606
rect 48837 298516 48865 298544
rect 48899 298516 48927 298544
rect 48961 298516 48989 298544
rect 49023 298516 49051 298544
rect 48837 298454 48865 298482
rect 48899 298454 48927 298482
rect 48961 298454 48989 298482
rect 49023 298454 49051 298482
rect 48837 298392 48865 298420
rect 48899 298392 48927 298420
rect 48961 298392 48989 298420
rect 49023 298392 49051 298420
rect 48837 290147 48865 290175
rect 48899 290147 48927 290175
rect 48961 290147 48989 290175
rect 49023 290147 49051 290175
rect 48837 290085 48865 290113
rect 48899 290085 48927 290113
rect 48961 290085 48989 290113
rect 49023 290085 49051 290113
rect 48837 290023 48865 290051
rect 48899 290023 48927 290051
rect 48961 290023 48989 290051
rect 49023 290023 49051 290051
rect 48837 289961 48865 289989
rect 48899 289961 48927 289989
rect 48961 289961 48989 289989
rect 49023 289961 49051 289989
rect 48837 281147 48865 281175
rect 48899 281147 48927 281175
rect 48961 281147 48989 281175
rect 49023 281147 49051 281175
rect 48837 281085 48865 281113
rect 48899 281085 48927 281113
rect 48961 281085 48989 281113
rect 49023 281085 49051 281113
rect 48837 281023 48865 281051
rect 48899 281023 48927 281051
rect 48961 281023 48989 281051
rect 49023 281023 49051 281051
rect 48837 280961 48865 280989
rect 48899 280961 48927 280989
rect 48961 280961 48989 280989
rect 49023 280961 49051 280989
rect 48837 272147 48865 272175
rect 48899 272147 48927 272175
rect 48961 272147 48989 272175
rect 49023 272147 49051 272175
rect 48837 272085 48865 272113
rect 48899 272085 48927 272113
rect 48961 272085 48989 272113
rect 49023 272085 49051 272113
rect 48837 272023 48865 272051
rect 48899 272023 48927 272051
rect 48961 272023 48989 272051
rect 49023 272023 49051 272051
rect 48837 271961 48865 271989
rect 48899 271961 48927 271989
rect 48961 271961 48989 271989
rect 49023 271961 49051 271989
rect 48837 263147 48865 263175
rect 48899 263147 48927 263175
rect 48961 263147 48989 263175
rect 49023 263147 49051 263175
rect 48837 263085 48865 263113
rect 48899 263085 48927 263113
rect 48961 263085 48989 263113
rect 49023 263085 49051 263113
rect 48837 263023 48865 263051
rect 48899 263023 48927 263051
rect 48961 263023 48989 263051
rect 49023 263023 49051 263051
rect 48837 262961 48865 262989
rect 48899 262961 48927 262989
rect 48961 262961 48989 262989
rect 49023 262961 49051 262989
rect 48837 254147 48865 254175
rect 48899 254147 48927 254175
rect 48961 254147 48989 254175
rect 49023 254147 49051 254175
rect 48837 254085 48865 254113
rect 48899 254085 48927 254113
rect 48961 254085 48989 254113
rect 49023 254085 49051 254113
rect 48837 254023 48865 254051
rect 48899 254023 48927 254051
rect 48961 254023 48989 254051
rect 49023 254023 49051 254051
rect 48837 253961 48865 253989
rect 48899 253961 48927 253989
rect 48961 253961 48989 253989
rect 49023 253961 49051 253989
rect 48837 245147 48865 245175
rect 48899 245147 48927 245175
rect 48961 245147 48989 245175
rect 49023 245147 49051 245175
rect 48837 245085 48865 245113
rect 48899 245085 48927 245113
rect 48961 245085 48989 245113
rect 49023 245085 49051 245113
rect 48837 245023 48865 245051
rect 48899 245023 48927 245051
rect 48961 245023 48989 245051
rect 49023 245023 49051 245051
rect 48837 244961 48865 244989
rect 48899 244961 48927 244989
rect 48961 244961 48989 244989
rect 49023 244961 49051 244989
rect 48837 236147 48865 236175
rect 48899 236147 48927 236175
rect 48961 236147 48989 236175
rect 49023 236147 49051 236175
rect 48837 236085 48865 236113
rect 48899 236085 48927 236113
rect 48961 236085 48989 236113
rect 49023 236085 49051 236113
rect 48837 236023 48865 236051
rect 48899 236023 48927 236051
rect 48961 236023 48989 236051
rect 49023 236023 49051 236051
rect 48837 235961 48865 235989
rect 48899 235961 48927 235989
rect 48961 235961 48989 235989
rect 49023 235961 49051 235989
rect 48837 227147 48865 227175
rect 48899 227147 48927 227175
rect 48961 227147 48989 227175
rect 49023 227147 49051 227175
rect 48837 227085 48865 227113
rect 48899 227085 48927 227113
rect 48961 227085 48989 227113
rect 49023 227085 49051 227113
rect 48837 227023 48865 227051
rect 48899 227023 48927 227051
rect 48961 227023 48989 227051
rect 49023 227023 49051 227051
rect 48837 226961 48865 226989
rect 48899 226961 48927 226989
rect 48961 226961 48989 226989
rect 49023 226961 49051 226989
rect 48837 218147 48865 218175
rect 48899 218147 48927 218175
rect 48961 218147 48989 218175
rect 49023 218147 49051 218175
rect 48837 218085 48865 218113
rect 48899 218085 48927 218113
rect 48961 218085 48989 218113
rect 49023 218085 49051 218113
rect 48837 218023 48865 218051
rect 48899 218023 48927 218051
rect 48961 218023 48989 218051
rect 49023 218023 49051 218051
rect 48837 217961 48865 217989
rect 48899 217961 48927 217989
rect 48961 217961 48989 217989
rect 49023 217961 49051 217989
rect 48837 209147 48865 209175
rect 48899 209147 48927 209175
rect 48961 209147 48989 209175
rect 49023 209147 49051 209175
rect 48837 209085 48865 209113
rect 48899 209085 48927 209113
rect 48961 209085 48989 209113
rect 49023 209085 49051 209113
rect 48837 209023 48865 209051
rect 48899 209023 48927 209051
rect 48961 209023 48989 209051
rect 49023 209023 49051 209051
rect 48837 208961 48865 208989
rect 48899 208961 48927 208989
rect 48961 208961 48989 208989
rect 49023 208961 49051 208989
rect 48837 200147 48865 200175
rect 48899 200147 48927 200175
rect 48961 200147 48989 200175
rect 49023 200147 49051 200175
rect 48837 200085 48865 200113
rect 48899 200085 48927 200113
rect 48961 200085 48989 200113
rect 49023 200085 49051 200113
rect 48837 200023 48865 200051
rect 48899 200023 48927 200051
rect 48961 200023 48989 200051
rect 49023 200023 49051 200051
rect 48837 199961 48865 199989
rect 48899 199961 48927 199989
rect 48961 199961 48989 199989
rect 49023 199961 49051 199989
rect 48837 191147 48865 191175
rect 48899 191147 48927 191175
rect 48961 191147 48989 191175
rect 49023 191147 49051 191175
rect 48837 191085 48865 191113
rect 48899 191085 48927 191113
rect 48961 191085 48989 191113
rect 49023 191085 49051 191113
rect 48837 191023 48865 191051
rect 48899 191023 48927 191051
rect 48961 191023 48989 191051
rect 49023 191023 49051 191051
rect 48837 190961 48865 190989
rect 48899 190961 48927 190989
rect 48961 190961 48989 190989
rect 49023 190961 49051 190989
rect 48837 182147 48865 182175
rect 48899 182147 48927 182175
rect 48961 182147 48989 182175
rect 49023 182147 49051 182175
rect 48837 182085 48865 182113
rect 48899 182085 48927 182113
rect 48961 182085 48989 182113
rect 49023 182085 49051 182113
rect 48837 182023 48865 182051
rect 48899 182023 48927 182051
rect 48961 182023 48989 182051
rect 49023 182023 49051 182051
rect 48837 181961 48865 181989
rect 48899 181961 48927 181989
rect 48961 181961 48989 181989
rect 49023 181961 49051 181989
rect 48837 173147 48865 173175
rect 48899 173147 48927 173175
rect 48961 173147 48989 173175
rect 49023 173147 49051 173175
rect 48837 173085 48865 173113
rect 48899 173085 48927 173113
rect 48961 173085 48989 173113
rect 49023 173085 49051 173113
rect 48837 173023 48865 173051
rect 48899 173023 48927 173051
rect 48961 173023 48989 173051
rect 49023 173023 49051 173051
rect 48837 172961 48865 172989
rect 48899 172961 48927 172989
rect 48961 172961 48989 172989
rect 49023 172961 49051 172989
rect 48837 164147 48865 164175
rect 48899 164147 48927 164175
rect 48961 164147 48989 164175
rect 49023 164147 49051 164175
rect 48837 164085 48865 164113
rect 48899 164085 48927 164113
rect 48961 164085 48989 164113
rect 49023 164085 49051 164113
rect 48837 164023 48865 164051
rect 48899 164023 48927 164051
rect 48961 164023 48989 164051
rect 49023 164023 49051 164051
rect 48837 163961 48865 163989
rect 48899 163961 48927 163989
rect 48961 163961 48989 163989
rect 49023 163961 49051 163989
rect 48837 155147 48865 155175
rect 48899 155147 48927 155175
rect 48961 155147 48989 155175
rect 49023 155147 49051 155175
rect 48837 155085 48865 155113
rect 48899 155085 48927 155113
rect 48961 155085 48989 155113
rect 49023 155085 49051 155113
rect 48837 155023 48865 155051
rect 48899 155023 48927 155051
rect 48961 155023 48989 155051
rect 49023 155023 49051 155051
rect 48837 154961 48865 154989
rect 48899 154961 48927 154989
rect 48961 154961 48989 154989
rect 49023 154961 49051 154989
rect 48837 146147 48865 146175
rect 48899 146147 48927 146175
rect 48961 146147 48989 146175
rect 49023 146147 49051 146175
rect 48837 146085 48865 146113
rect 48899 146085 48927 146113
rect 48961 146085 48989 146113
rect 49023 146085 49051 146113
rect 48837 146023 48865 146051
rect 48899 146023 48927 146051
rect 48961 146023 48989 146051
rect 49023 146023 49051 146051
rect 48837 145961 48865 145989
rect 48899 145961 48927 145989
rect 48961 145961 48989 145989
rect 49023 145961 49051 145989
rect 48837 137147 48865 137175
rect 48899 137147 48927 137175
rect 48961 137147 48989 137175
rect 49023 137147 49051 137175
rect 48837 137085 48865 137113
rect 48899 137085 48927 137113
rect 48961 137085 48989 137113
rect 49023 137085 49051 137113
rect 48837 137023 48865 137051
rect 48899 137023 48927 137051
rect 48961 137023 48989 137051
rect 49023 137023 49051 137051
rect 48837 136961 48865 136989
rect 48899 136961 48927 136989
rect 48961 136961 48989 136989
rect 49023 136961 49051 136989
rect 48837 128147 48865 128175
rect 48899 128147 48927 128175
rect 48961 128147 48989 128175
rect 49023 128147 49051 128175
rect 48837 128085 48865 128113
rect 48899 128085 48927 128113
rect 48961 128085 48989 128113
rect 49023 128085 49051 128113
rect 48837 128023 48865 128051
rect 48899 128023 48927 128051
rect 48961 128023 48989 128051
rect 49023 128023 49051 128051
rect 48837 127961 48865 127989
rect 48899 127961 48927 127989
rect 48961 127961 48989 127989
rect 49023 127961 49051 127989
rect 48837 119147 48865 119175
rect 48899 119147 48927 119175
rect 48961 119147 48989 119175
rect 49023 119147 49051 119175
rect 48837 119085 48865 119113
rect 48899 119085 48927 119113
rect 48961 119085 48989 119113
rect 49023 119085 49051 119113
rect 48837 119023 48865 119051
rect 48899 119023 48927 119051
rect 48961 119023 48989 119051
rect 49023 119023 49051 119051
rect 48837 118961 48865 118989
rect 48899 118961 48927 118989
rect 48961 118961 48989 118989
rect 49023 118961 49051 118989
rect 48837 110147 48865 110175
rect 48899 110147 48927 110175
rect 48961 110147 48989 110175
rect 49023 110147 49051 110175
rect 48837 110085 48865 110113
rect 48899 110085 48927 110113
rect 48961 110085 48989 110113
rect 49023 110085 49051 110113
rect 48837 110023 48865 110051
rect 48899 110023 48927 110051
rect 48961 110023 48989 110051
rect 49023 110023 49051 110051
rect 48837 109961 48865 109989
rect 48899 109961 48927 109989
rect 48961 109961 48989 109989
rect 49023 109961 49051 109989
rect 48837 101147 48865 101175
rect 48899 101147 48927 101175
rect 48961 101147 48989 101175
rect 49023 101147 49051 101175
rect 48837 101085 48865 101113
rect 48899 101085 48927 101113
rect 48961 101085 48989 101113
rect 49023 101085 49051 101113
rect 48837 101023 48865 101051
rect 48899 101023 48927 101051
rect 48961 101023 48989 101051
rect 49023 101023 49051 101051
rect 48837 100961 48865 100989
rect 48899 100961 48927 100989
rect 48961 100961 48989 100989
rect 49023 100961 49051 100989
rect 48837 92147 48865 92175
rect 48899 92147 48927 92175
rect 48961 92147 48989 92175
rect 49023 92147 49051 92175
rect 48837 92085 48865 92113
rect 48899 92085 48927 92113
rect 48961 92085 48989 92113
rect 49023 92085 49051 92113
rect 48837 92023 48865 92051
rect 48899 92023 48927 92051
rect 48961 92023 48989 92051
rect 49023 92023 49051 92051
rect 48837 91961 48865 91989
rect 48899 91961 48927 91989
rect 48961 91961 48989 91989
rect 49023 91961 49051 91989
rect 48837 83147 48865 83175
rect 48899 83147 48927 83175
rect 48961 83147 48989 83175
rect 49023 83147 49051 83175
rect 48837 83085 48865 83113
rect 48899 83085 48927 83113
rect 48961 83085 48989 83113
rect 49023 83085 49051 83113
rect 48837 83023 48865 83051
rect 48899 83023 48927 83051
rect 48961 83023 48989 83051
rect 49023 83023 49051 83051
rect 48837 82961 48865 82989
rect 48899 82961 48927 82989
rect 48961 82961 48989 82989
rect 49023 82961 49051 82989
rect 48837 74147 48865 74175
rect 48899 74147 48927 74175
rect 48961 74147 48989 74175
rect 49023 74147 49051 74175
rect 48837 74085 48865 74113
rect 48899 74085 48927 74113
rect 48961 74085 48989 74113
rect 49023 74085 49051 74113
rect 48837 74023 48865 74051
rect 48899 74023 48927 74051
rect 48961 74023 48989 74051
rect 49023 74023 49051 74051
rect 48837 73961 48865 73989
rect 48899 73961 48927 73989
rect 48961 73961 48989 73989
rect 49023 73961 49051 73989
rect 48837 65147 48865 65175
rect 48899 65147 48927 65175
rect 48961 65147 48989 65175
rect 49023 65147 49051 65175
rect 48837 65085 48865 65113
rect 48899 65085 48927 65113
rect 48961 65085 48989 65113
rect 49023 65085 49051 65113
rect 48837 65023 48865 65051
rect 48899 65023 48927 65051
rect 48961 65023 48989 65051
rect 49023 65023 49051 65051
rect 48837 64961 48865 64989
rect 48899 64961 48927 64989
rect 48961 64961 48989 64989
rect 49023 64961 49051 64989
rect 48837 56147 48865 56175
rect 48899 56147 48927 56175
rect 48961 56147 48989 56175
rect 49023 56147 49051 56175
rect 48837 56085 48865 56113
rect 48899 56085 48927 56113
rect 48961 56085 48989 56113
rect 49023 56085 49051 56113
rect 48837 56023 48865 56051
rect 48899 56023 48927 56051
rect 48961 56023 48989 56051
rect 49023 56023 49051 56051
rect 48837 55961 48865 55989
rect 48899 55961 48927 55989
rect 48961 55961 48989 55989
rect 49023 55961 49051 55989
rect 48837 47147 48865 47175
rect 48899 47147 48927 47175
rect 48961 47147 48989 47175
rect 49023 47147 49051 47175
rect 48837 47085 48865 47113
rect 48899 47085 48927 47113
rect 48961 47085 48989 47113
rect 49023 47085 49051 47113
rect 48837 47023 48865 47051
rect 48899 47023 48927 47051
rect 48961 47023 48989 47051
rect 49023 47023 49051 47051
rect 48837 46961 48865 46989
rect 48899 46961 48927 46989
rect 48961 46961 48989 46989
rect 49023 46961 49051 46989
rect 48837 38147 48865 38175
rect 48899 38147 48927 38175
rect 48961 38147 48989 38175
rect 49023 38147 49051 38175
rect 48837 38085 48865 38113
rect 48899 38085 48927 38113
rect 48961 38085 48989 38113
rect 49023 38085 49051 38113
rect 48837 38023 48865 38051
rect 48899 38023 48927 38051
rect 48961 38023 48989 38051
rect 49023 38023 49051 38051
rect 48837 37961 48865 37989
rect 48899 37961 48927 37989
rect 48961 37961 48989 37989
rect 49023 37961 49051 37989
rect 48837 29147 48865 29175
rect 48899 29147 48927 29175
rect 48961 29147 48989 29175
rect 49023 29147 49051 29175
rect 48837 29085 48865 29113
rect 48899 29085 48927 29113
rect 48961 29085 48989 29113
rect 49023 29085 49051 29113
rect 48837 29023 48865 29051
rect 48899 29023 48927 29051
rect 48961 29023 48989 29051
rect 49023 29023 49051 29051
rect 48837 28961 48865 28989
rect 48899 28961 48927 28989
rect 48961 28961 48989 28989
rect 49023 28961 49051 28989
rect 48837 20147 48865 20175
rect 48899 20147 48927 20175
rect 48961 20147 48989 20175
rect 49023 20147 49051 20175
rect 48837 20085 48865 20113
rect 48899 20085 48927 20113
rect 48961 20085 48989 20113
rect 49023 20085 49051 20113
rect 48837 20023 48865 20051
rect 48899 20023 48927 20051
rect 48961 20023 48989 20051
rect 49023 20023 49051 20051
rect 48837 19961 48865 19989
rect 48899 19961 48927 19989
rect 48961 19961 48989 19989
rect 49023 19961 49051 19989
rect 48837 11147 48865 11175
rect 48899 11147 48927 11175
rect 48961 11147 48989 11175
rect 49023 11147 49051 11175
rect 48837 11085 48865 11113
rect 48899 11085 48927 11113
rect 48961 11085 48989 11113
rect 49023 11085 49051 11113
rect 48837 11023 48865 11051
rect 48899 11023 48927 11051
rect 48961 11023 48989 11051
rect 49023 11023 49051 11051
rect 48837 10961 48865 10989
rect 48899 10961 48927 10989
rect 48961 10961 48989 10989
rect 49023 10961 49051 10989
rect 48837 2147 48865 2175
rect 48899 2147 48927 2175
rect 48961 2147 48989 2175
rect 49023 2147 49051 2175
rect 48837 2085 48865 2113
rect 48899 2085 48927 2113
rect 48961 2085 48989 2113
rect 49023 2085 49051 2113
rect 48837 2023 48865 2051
rect 48899 2023 48927 2051
rect 48961 2023 48989 2051
rect 49023 2023 49051 2051
rect 48837 1961 48865 1989
rect 48899 1961 48927 1989
rect 48961 1961 48989 1989
rect 49023 1961 49051 1989
rect 48837 -108 48865 -80
rect 48899 -108 48927 -80
rect 48961 -108 48989 -80
rect 49023 -108 49051 -80
rect 48837 -170 48865 -142
rect 48899 -170 48927 -142
rect 48961 -170 48989 -142
rect 49023 -170 49051 -142
rect 48837 -232 48865 -204
rect 48899 -232 48927 -204
rect 48961 -232 48989 -204
rect 49023 -232 49051 -204
rect 48837 -294 48865 -266
rect 48899 -294 48927 -266
rect 48961 -294 48989 -266
rect 49023 -294 49051 -266
rect 50697 299058 50725 299086
rect 50759 299058 50787 299086
rect 50821 299058 50849 299086
rect 50883 299058 50911 299086
rect 50697 298996 50725 299024
rect 50759 298996 50787 299024
rect 50821 298996 50849 299024
rect 50883 298996 50911 299024
rect 50697 298934 50725 298962
rect 50759 298934 50787 298962
rect 50821 298934 50849 298962
rect 50883 298934 50911 298962
rect 50697 298872 50725 298900
rect 50759 298872 50787 298900
rect 50821 298872 50849 298900
rect 50883 298872 50911 298900
rect 50697 293147 50725 293175
rect 50759 293147 50787 293175
rect 50821 293147 50849 293175
rect 50883 293147 50911 293175
rect 50697 293085 50725 293113
rect 50759 293085 50787 293113
rect 50821 293085 50849 293113
rect 50883 293085 50911 293113
rect 50697 293023 50725 293051
rect 50759 293023 50787 293051
rect 50821 293023 50849 293051
rect 50883 293023 50911 293051
rect 50697 292961 50725 292989
rect 50759 292961 50787 292989
rect 50821 292961 50849 292989
rect 50883 292961 50911 292989
rect 50697 284147 50725 284175
rect 50759 284147 50787 284175
rect 50821 284147 50849 284175
rect 50883 284147 50911 284175
rect 50697 284085 50725 284113
rect 50759 284085 50787 284113
rect 50821 284085 50849 284113
rect 50883 284085 50911 284113
rect 50697 284023 50725 284051
rect 50759 284023 50787 284051
rect 50821 284023 50849 284051
rect 50883 284023 50911 284051
rect 50697 283961 50725 283989
rect 50759 283961 50787 283989
rect 50821 283961 50849 283989
rect 50883 283961 50911 283989
rect 50697 275147 50725 275175
rect 50759 275147 50787 275175
rect 50821 275147 50849 275175
rect 50883 275147 50911 275175
rect 50697 275085 50725 275113
rect 50759 275085 50787 275113
rect 50821 275085 50849 275113
rect 50883 275085 50911 275113
rect 50697 275023 50725 275051
rect 50759 275023 50787 275051
rect 50821 275023 50849 275051
rect 50883 275023 50911 275051
rect 50697 274961 50725 274989
rect 50759 274961 50787 274989
rect 50821 274961 50849 274989
rect 50883 274961 50911 274989
rect 50697 266147 50725 266175
rect 50759 266147 50787 266175
rect 50821 266147 50849 266175
rect 50883 266147 50911 266175
rect 50697 266085 50725 266113
rect 50759 266085 50787 266113
rect 50821 266085 50849 266113
rect 50883 266085 50911 266113
rect 50697 266023 50725 266051
rect 50759 266023 50787 266051
rect 50821 266023 50849 266051
rect 50883 266023 50911 266051
rect 50697 265961 50725 265989
rect 50759 265961 50787 265989
rect 50821 265961 50849 265989
rect 50883 265961 50911 265989
rect 50697 257147 50725 257175
rect 50759 257147 50787 257175
rect 50821 257147 50849 257175
rect 50883 257147 50911 257175
rect 50697 257085 50725 257113
rect 50759 257085 50787 257113
rect 50821 257085 50849 257113
rect 50883 257085 50911 257113
rect 50697 257023 50725 257051
rect 50759 257023 50787 257051
rect 50821 257023 50849 257051
rect 50883 257023 50911 257051
rect 50697 256961 50725 256989
rect 50759 256961 50787 256989
rect 50821 256961 50849 256989
rect 50883 256961 50911 256989
rect 50697 248147 50725 248175
rect 50759 248147 50787 248175
rect 50821 248147 50849 248175
rect 50883 248147 50911 248175
rect 50697 248085 50725 248113
rect 50759 248085 50787 248113
rect 50821 248085 50849 248113
rect 50883 248085 50911 248113
rect 50697 248023 50725 248051
rect 50759 248023 50787 248051
rect 50821 248023 50849 248051
rect 50883 248023 50911 248051
rect 50697 247961 50725 247989
rect 50759 247961 50787 247989
rect 50821 247961 50849 247989
rect 50883 247961 50911 247989
rect 50697 239147 50725 239175
rect 50759 239147 50787 239175
rect 50821 239147 50849 239175
rect 50883 239147 50911 239175
rect 50697 239085 50725 239113
rect 50759 239085 50787 239113
rect 50821 239085 50849 239113
rect 50883 239085 50911 239113
rect 50697 239023 50725 239051
rect 50759 239023 50787 239051
rect 50821 239023 50849 239051
rect 50883 239023 50911 239051
rect 50697 238961 50725 238989
rect 50759 238961 50787 238989
rect 50821 238961 50849 238989
rect 50883 238961 50911 238989
rect 50697 230147 50725 230175
rect 50759 230147 50787 230175
rect 50821 230147 50849 230175
rect 50883 230147 50911 230175
rect 50697 230085 50725 230113
rect 50759 230085 50787 230113
rect 50821 230085 50849 230113
rect 50883 230085 50911 230113
rect 50697 230023 50725 230051
rect 50759 230023 50787 230051
rect 50821 230023 50849 230051
rect 50883 230023 50911 230051
rect 50697 229961 50725 229989
rect 50759 229961 50787 229989
rect 50821 229961 50849 229989
rect 50883 229961 50911 229989
rect 50697 221147 50725 221175
rect 50759 221147 50787 221175
rect 50821 221147 50849 221175
rect 50883 221147 50911 221175
rect 50697 221085 50725 221113
rect 50759 221085 50787 221113
rect 50821 221085 50849 221113
rect 50883 221085 50911 221113
rect 50697 221023 50725 221051
rect 50759 221023 50787 221051
rect 50821 221023 50849 221051
rect 50883 221023 50911 221051
rect 50697 220961 50725 220989
rect 50759 220961 50787 220989
rect 50821 220961 50849 220989
rect 50883 220961 50911 220989
rect 50697 212147 50725 212175
rect 50759 212147 50787 212175
rect 50821 212147 50849 212175
rect 50883 212147 50911 212175
rect 50697 212085 50725 212113
rect 50759 212085 50787 212113
rect 50821 212085 50849 212113
rect 50883 212085 50911 212113
rect 50697 212023 50725 212051
rect 50759 212023 50787 212051
rect 50821 212023 50849 212051
rect 50883 212023 50911 212051
rect 50697 211961 50725 211989
rect 50759 211961 50787 211989
rect 50821 211961 50849 211989
rect 50883 211961 50911 211989
rect 50697 203147 50725 203175
rect 50759 203147 50787 203175
rect 50821 203147 50849 203175
rect 50883 203147 50911 203175
rect 50697 203085 50725 203113
rect 50759 203085 50787 203113
rect 50821 203085 50849 203113
rect 50883 203085 50911 203113
rect 50697 203023 50725 203051
rect 50759 203023 50787 203051
rect 50821 203023 50849 203051
rect 50883 203023 50911 203051
rect 50697 202961 50725 202989
rect 50759 202961 50787 202989
rect 50821 202961 50849 202989
rect 50883 202961 50911 202989
rect 50697 194147 50725 194175
rect 50759 194147 50787 194175
rect 50821 194147 50849 194175
rect 50883 194147 50911 194175
rect 50697 194085 50725 194113
rect 50759 194085 50787 194113
rect 50821 194085 50849 194113
rect 50883 194085 50911 194113
rect 50697 194023 50725 194051
rect 50759 194023 50787 194051
rect 50821 194023 50849 194051
rect 50883 194023 50911 194051
rect 50697 193961 50725 193989
rect 50759 193961 50787 193989
rect 50821 193961 50849 193989
rect 50883 193961 50911 193989
rect 50697 185147 50725 185175
rect 50759 185147 50787 185175
rect 50821 185147 50849 185175
rect 50883 185147 50911 185175
rect 50697 185085 50725 185113
rect 50759 185085 50787 185113
rect 50821 185085 50849 185113
rect 50883 185085 50911 185113
rect 50697 185023 50725 185051
rect 50759 185023 50787 185051
rect 50821 185023 50849 185051
rect 50883 185023 50911 185051
rect 50697 184961 50725 184989
rect 50759 184961 50787 184989
rect 50821 184961 50849 184989
rect 50883 184961 50911 184989
rect 50697 176147 50725 176175
rect 50759 176147 50787 176175
rect 50821 176147 50849 176175
rect 50883 176147 50911 176175
rect 50697 176085 50725 176113
rect 50759 176085 50787 176113
rect 50821 176085 50849 176113
rect 50883 176085 50911 176113
rect 50697 176023 50725 176051
rect 50759 176023 50787 176051
rect 50821 176023 50849 176051
rect 50883 176023 50911 176051
rect 50697 175961 50725 175989
rect 50759 175961 50787 175989
rect 50821 175961 50849 175989
rect 50883 175961 50911 175989
rect 50697 167147 50725 167175
rect 50759 167147 50787 167175
rect 50821 167147 50849 167175
rect 50883 167147 50911 167175
rect 50697 167085 50725 167113
rect 50759 167085 50787 167113
rect 50821 167085 50849 167113
rect 50883 167085 50911 167113
rect 50697 167023 50725 167051
rect 50759 167023 50787 167051
rect 50821 167023 50849 167051
rect 50883 167023 50911 167051
rect 50697 166961 50725 166989
rect 50759 166961 50787 166989
rect 50821 166961 50849 166989
rect 50883 166961 50911 166989
rect 50697 158147 50725 158175
rect 50759 158147 50787 158175
rect 50821 158147 50849 158175
rect 50883 158147 50911 158175
rect 50697 158085 50725 158113
rect 50759 158085 50787 158113
rect 50821 158085 50849 158113
rect 50883 158085 50911 158113
rect 50697 158023 50725 158051
rect 50759 158023 50787 158051
rect 50821 158023 50849 158051
rect 50883 158023 50911 158051
rect 50697 157961 50725 157989
rect 50759 157961 50787 157989
rect 50821 157961 50849 157989
rect 50883 157961 50911 157989
rect 50697 149147 50725 149175
rect 50759 149147 50787 149175
rect 50821 149147 50849 149175
rect 50883 149147 50911 149175
rect 50697 149085 50725 149113
rect 50759 149085 50787 149113
rect 50821 149085 50849 149113
rect 50883 149085 50911 149113
rect 50697 149023 50725 149051
rect 50759 149023 50787 149051
rect 50821 149023 50849 149051
rect 50883 149023 50911 149051
rect 50697 148961 50725 148989
rect 50759 148961 50787 148989
rect 50821 148961 50849 148989
rect 50883 148961 50911 148989
rect 50697 140147 50725 140175
rect 50759 140147 50787 140175
rect 50821 140147 50849 140175
rect 50883 140147 50911 140175
rect 50697 140085 50725 140113
rect 50759 140085 50787 140113
rect 50821 140085 50849 140113
rect 50883 140085 50911 140113
rect 50697 140023 50725 140051
rect 50759 140023 50787 140051
rect 50821 140023 50849 140051
rect 50883 140023 50911 140051
rect 50697 139961 50725 139989
rect 50759 139961 50787 139989
rect 50821 139961 50849 139989
rect 50883 139961 50911 139989
rect 50697 131147 50725 131175
rect 50759 131147 50787 131175
rect 50821 131147 50849 131175
rect 50883 131147 50911 131175
rect 50697 131085 50725 131113
rect 50759 131085 50787 131113
rect 50821 131085 50849 131113
rect 50883 131085 50911 131113
rect 50697 131023 50725 131051
rect 50759 131023 50787 131051
rect 50821 131023 50849 131051
rect 50883 131023 50911 131051
rect 50697 130961 50725 130989
rect 50759 130961 50787 130989
rect 50821 130961 50849 130989
rect 50883 130961 50911 130989
rect 50697 122147 50725 122175
rect 50759 122147 50787 122175
rect 50821 122147 50849 122175
rect 50883 122147 50911 122175
rect 50697 122085 50725 122113
rect 50759 122085 50787 122113
rect 50821 122085 50849 122113
rect 50883 122085 50911 122113
rect 50697 122023 50725 122051
rect 50759 122023 50787 122051
rect 50821 122023 50849 122051
rect 50883 122023 50911 122051
rect 50697 121961 50725 121989
rect 50759 121961 50787 121989
rect 50821 121961 50849 121989
rect 50883 121961 50911 121989
rect 50697 113147 50725 113175
rect 50759 113147 50787 113175
rect 50821 113147 50849 113175
rect 50883 113147 50911 113175
rect 50697 113085 50725 113113
rect 50759 113085 50787 113113
rect 50821 113085 50849 113113
rect 50883 113085 50911 113113
rect 50697 113023 50725 113051
rect 50759 113023 50787 113051
rect 50821 113023 50849 113051
rect 50883 113023 50911 113051
rect 50697 112961 50725 112989
rect 50759 112961 50787 112989
rect 50821 112961 50849 112989
rect 50883 112961 50911 112989
rect 50697 104147 50725 104175
rect 50759 104147 50787 104175
rect 50821 104147 50849 104175
rect 50883 104147 50911 104175
rect 50697 104085 50725 104113
rect 50759 104085 50787 104113
rect 50821 104085 50849 104113
rect 50883 104085 50911 104113
rect 50697 104023 50725 104051
rect 50759 104023 50787 104051
rect 50821 104023 50849 104051
rect 50883 104023 50911 104051
rect 50697 103961 50725 103989
rect 50759 103961 50787 103989
rect 50821 103961 50849 103989
rect 50883 103961 50911 103989
rect 50697 95147 50725 95175
rect 50759 95147 50787 95175
rect 50821 95147 50849 95175
rect 50883 95147 50911 95175
rect 50697 95085 50725 95113
rect 50759 95085 50787 95113
rect 50821 95085 50849 95113
rect 50883 95085 50911 95113
rect 50697 95023 50725 95051
rect 50759 95023 50787 95051
rect 50821 95023 50849 95051
rect 50883 95023 50911 95051
rect 50697 94961 50725 94989
rect 50759 94961 50787 94989
rect 50821 94961 50849 94989
rect 50883 94961 50911 94989
rect 50697 86147 50725 86175
rect 50759 86147 50787 86175
rect 50821 86147 50849 86175
rect 50883 86147 50911 86175
rect 50697 86085 50725 86113
rect 50759 86085 50787 86113
rect 50821 86085 50849 86113
rect 50883 86085 50911 86113
rect 50697 86023 50725 86051
rect 50759 86023 50787 86051
rect 50821 86023 50849 86051
rect 50883 86023 50911 86051
rect 50697 85961 50725 85989
rect 50759 85961 50787 85989
rect 50821 85961 50849 85989
rect 50883 85961 50911 85989
rect 50697 77147 50725 77175
rect 50759 77147 50787 77175
rect 50821 77147 50849 77175
rect 50883 77147 50911 77175
rect 50697 77085 50725 77113
rect 50759 77085 50787 77113
rect 50821 77085 50849 77113
rect 50883 77085 50911 77113
rect 50697 77023 50725 77051
rect 50759 77023 50787 77051
rect 50821 77023 50849 77051
rect 50883 77023 50911 77051
rect 50697 76961 50725 76989
rect 50759 76961 50787 76989
rect 50821 76961 50849 76989
rect 50883 76961 50911 76989
rect 50697 68147 50725 68175
rect 50759 68147 50787 68175
rect 50821 68147 50849 68175
rect 50883 68147 50911 68175
rect 50697 68085 50725 68113
rect 50759 68085 50787 68113
rect 50821 68085 50849 68113
rect 50883 68085 50911 68113
rect 50697 68023 50725 68051
rect 50759 68023 50787 68051
rect 50821 68023 50849 68051
rect 50883 68023 50911 68051
rect 50697 67961 50725 67989
rect 50759 67961 50787 67989
rect 50821 67961 50849 67989
rect 50883 67961 50911 67989
rect 50697 59147 50725 59175
rect 50759 59147 50787 59175
rect 50821 59147 50849 59175
rect 50883 59147 50911 59175
rect 50697 59085 50725 59113
rect 50759 59085 50787 59113
rect 50821 59085 50849 59113
rect 50883 59085 50911 59113
rect 50697 59023 50725 59051
rect 50759 59023 50787 59051
rect 50821 59023 50849 59051
rect 50883 59023 50911 59051
rect 50697 58961 50725 58989
rect 50759 58961 50787 58989
rect 50821 58961 50849 58989
rect 50883 58961 50911 58989
rect 50697 50147 50725 50175
rect 50759 50147 50787 50175
rect 50821 50147 50849 50175
rect 50883 50147 50911 50175
rect 50697 50085 50725 50113
rect 50759 50085 50787 50113
rect 50821 50085 50849 50113
rect 50883 50085 50911 50113
rect 50697 50023 50725 50051
rect 50759 50023 50787 50051
rect 50821 50023 50849 50051
rect 50883 50023 50911 50051
rect 50697 49961 50725 49989
rect 50759 49961 50787 49989
rect 50821 49961 50849 49989
rect 50883 49961 50911 49989
rect 50697 41147 50725 41175
rect 50759 41147 50787 41175
rect 50821 41147 50849 41175
rect 50883 41147 50911 41175
rect 50697 41085 50725 41113
rect 50759 41085 50787 41113
rect 50821 41085 50849 41113
rect 50883 41085 50911 41113
rect 50697 41023 50725 41051
rect 50759 41023 50787 41051
rect 50821 41023 50849 41051
rect 50883 41023 50911 41051
rect 50697 40961 50725 40989
rect 50759 40961 50787 40989
rect 50821 40961 50849 40989
rect 50883 40961 50911 40989
rect 50697 32147 50725 32175
rect 50759 32147 50787 32175
rect 50821 32147 50849 32175
rect 50883 32147 50911 32175
rect 50697 32085 50725 32113
rect 50759 32085 50787 32113
rect 50821 32085 50849 32113
rect 50883 32085 50911 32113
rect 50697 32023 50725 32051
rect 50759 32023 50787 32051
rect 50821 32023 50849 32051
rect 50883 32023 50911 32051
rect 50697 31961 50725 31989
rect 50759 31961 50787 31989
rect 50821 31961 50849 31989
rect 50883 31961 50911 31989
rect 50697 23147 50725 23175
rect 50759 23147 50787 23175
rect 50821 23147 50849 23175
rect 50883 23147 50911 23175
rect 50697 23085 50725 23113
rect 50759 23085 50787 23113
rect 50821 23085 50849 23113
rect 50883 23085 50911 23113
rect 50697 23023 50725 23051
rect 50759 23023 50787 23051
rect 50821 23023 50849 23051
rect 50883 23023 50911 23051
rect 50697 22961 50725 22989
rect 50759 22961 50787 22989
rect 50821 22961 50849 22989
rect 50883 22961 50911 22989
rect 50697 14147 50725 14175
rect 50759 14147 50787 14175
rect 50821 14147 50849 14175
rect 50883 14147 50911 14175
rect 50697 14085 50725 14113
rect 50759 14085 50787 14113
rect 50821 14085 50849 14113
rect 50883 14085 50911 14113
rect 50697 14023 50725 14051
rect 50759 14023 50787 14051
rect 50821 14023 50849 14051
rect 50883 14023 50911 14051
rect 50697 13961 50725 13989
rect 50759 13961 50787 13989
rect 50821 13961 50849 13989
rect 50883 13961 50911 13989
rect 50697 5147 50725 5175
rect 50759 5147 50787 5175
rect 50821 5147 50849 5175
rect 50883 5147 50911 5175
rect 50697 5085 50725 5113
rect 50759 5085 50787 5113
rect 50821 5085 50849 5113
rect 50883 5085 50911 5113
rect 50697 5023 50725 5051
rect 50759 5023 50787 5051
rect 50821 5023 50849 5051
rect 50883 5023 50911 5051
rect 50697 4961 50725 4989
rect 50759 4961 50787 4989
rect 50821 4961 50849 4989
rect 50883 4961 50911 4989
rect 50697 -588 50725 -560
rect 50759 -588 50787 -560
rect 50821 -588 50849 -560
rect 50883 -588 50911 -560
rect 50697 -650 50725 -622
rect 50759 -650 50787 -622
rect 50821 -650 50849 -622
rect 50883 -650 50911 -622
rect 50697 -712 50725 -684
rect 50759 -712 50787 -684
rect 50821 -712 50849 -684
rect 50883 -712 50911 -684
rect 50697 -774 50725 -746
rect 50759 -774 50787 -746
rect 50821 -774 50849 -746
rect 50883 -774 50911 -746
rect 64197 298578 64225 298606
rect 64259 298578 64287 298606
rect 64321 298578 64349 298606
rect 64383 298578 64411 298606
rect 64197 298516 64225 298544
rect 64259 298516 64287 298544
rect 64321 298516 64349 298544
rect 64383 298516 64411 298544
rect 64197 298454 64225 298482
rect 64259 298454 64287 298482
rect 64321 298454 64349 298482
rect 64383 298454 64411 298482
rect 64197 298392 64225 298420
rect 64259 298392 64287 298420
rect 64321 298392 64349 298420
rect 64383 298392 64411 298420
rect 64197 290147 64225 290175
rect 64259 290147 64287 290175
rect 64321 290147 64349 290175
rect 64383 290147 64411 290175
rect 64197 290085 64225 290113
rect 64259 290085 64287 290113
rect 64321 290085 64349 290113
rect 64383 290085 64411 290113
rect 64197 290023 64225 290051
rect 64259 290023 64287 290051
rect 64321 290023 64349 290051
rect 64383 290023 64411 290051
rect 64197 289961 64225 289989
rect 64259 289961 64287 289989
rect 64321 289961 64349 289989
rect 64383 289961 64411 289989
rect 64197 281147 64225 281175
rect 64259 281147 64287 281175
rect 64321 281147 64349 281175
rect 64383 281147 64411 281175
rect 64197 281085 64225 281113
rect 64259 281085 64287 281113
rect 64321 281085 64349 281113
rect 64383 281085 64411 281113
rect 64197 281023 64225 281051
rect 64259 281023 64287 281051
rect 64321 281023 64349 281051
rect 64383 281023 64411 281051
rect 64197 280961 64225 280989
rect 64259 280961 64287 280989
rect 64321 280961 64349 280989
rect 64383 280961 64411 280989
rect 64197 272147 64225 272175
rect 64259 272147 64287 272175
rect 64321 272147 64349 272175
rect 64383 272147 64411 272175
rect 64197 272085 64225 272113
rect 64259 272085 64287 272113
rect 64321 272085 64349 272113
rect 64383 272085 64411 272113
rect 64197 272023 64225 272051
rect 64259 272023 64287 272051
rect 64321 272023 64349 272051
rect 64383 272023 64411 272051
rect 64197 271961 64225 271989
rect 64259 271961 64287 271989
rect 64321 271961 64349 271989
rect 64383 271961 64411 271989
rect 64197 263147 64225 263175
rect 64259 263147 64287 263175
rect 64321 263147 64349 263175
rect 64383 263147 64411 263175
rect 64197 263085 64225 263113
rect 64259 263085 64287 263113
rect 64321 263085 64349 263113
rect 64383 263085 64411 263113
rect 64197 263023 64225 263051
rect 64259 263023 64287 263051
rect 64321 263023 64349 263051
rect 64383 263023 64411 263051
rect 64197 262961 64225 262989
rect 64259 262961 64287 262989
rect 64321 262961 64349 262989
rect 64383 262961 64411 262989
rect 64197 254147 64225 254175
rect 64259 254147 64287 254175
rect 64321 254147 64349 254175
rect 64383 254147 64411 254175
rect 64197 254085 64225 254113
rect 64259 254085 64287 254113
rect 64321 254085 64349 254113
rect 64383 254085 64411 254113
rect 64197 254023 64225 254051
rect 64259 254023 64287 254051
rect 64321 254023 64349 254051
rect 64383 254023 64411 254051
rect 64197 253961 64225 253989
rect 64259 253961 64287 253989
rect 64321 253961 64349 253989
rect 64383 253961 64411 253989
rect 64197 245147 64225 245175
rect 64259 245147 64287 245175
rect 64321 245147 64349 245175
rect 64383 245147 64411 245175
rect 64197 245085 64225 245113
rect 64259 245085 64287 245113
rect 64321 245085 64349 245113
rect 64383 245085 64411 245113
rect 64197 245023 64225 245051
rect 64259 245023 64287 245051
rect 64321 245023 64349 245051
rect 64383 245023 64411 245051
rect 64197 244961 64225 244989
rect 64259 244961 64287 244989
rect 64321 244961 64349 244989
rect 64383 244961 64411 244989
rect 64197 236147 64225 236175
rect 64259 236147 64287 236175
rect 64321 236147 64349 236175
rect 64383 236147 64411 236175
rect 64197 236085 64225 236113
rect 64259 236085 64287 236113
rect 64321 236085 64349 236113
rect 64383 236085 64411 236113
rect 64197 236023 64225 236051
rect 64259 236023 64287 236051
rect 64321 236023 64349 236051
rect 64383 236023 64411 236051
rect 64197 235961 64225 235989
rect 64259 235961 64287 235989
rect 64321 235961 64349 235989
rect 64383 235961 64411 235989
rect 64197 227147 64225 227175
rect 64259 227147 64287 227175
rect 64321 227147 64349 227175
rect 64383 227147 64411 227175
rect 64197 227085 64225 227113
rect 64259 227085 64287 227113
rect 64321 227085 64349 227113
rect 64383 227085 64411 227113
rect 64197 227023 64225 227051
rect 64259 227023 64287 227051
rect 64321 227023 64349 227051
rect 64383 227023 64411 227051
rect 64197 226961 64225 226989
rect 64259 226961 64287 226989
rect 64321 226961 64349 226989
rect 64383 226961 64411 226989
rect 64197 218147 64225 218175
rect 64259 218147 64287 218175
rect 64321 218147 64349 218175
rect 64383 218147 64411 218175
rect 64197 218085 64225 218113
rect 64259 218085 64287 218113
rect 64321 218085 64349 218113
rect 64383 218085 64411 218113
rect 64197 218023 64225 218051
rect 64259 218023 64287 218051
rect 64321 218023 64349 218051
rect 64383 218023 64411 218051
rect 64197 217961 64225 217989
rect 64259 217961 64287 217989
rect 64321 217961 64349 217989
rect 64383 217961 64411 217989
rect 64197 209147 64225 209175
rect 64259 209147 64287 209175
rect 64321 209147 64349 209175
rect 64383 209147 64411 209175
rect 64197 209085 64225 209113
rect 64259 209085 64287 209113
rect 64321 209085 64349 209113
rect 64383 209085 64411 209113
rect 64197 209023 64225 209051
rect 64259 209023 64287 209051
rect 64321 209023 64349 209051
rect 64383 209023 64411 209051
rect 64197 208961 64225 208989
rect 64259 208961 64287 208989
rect 64321 208961 64349 208989
rect 64383 208961 64411 208989
rect 64197 200147 64225 200175
rect 64259 200147 64287 200175
rect 64321 200147 64349 200175
rect 64383 200147 64411 200175
rect 64197 200085 64225 200113
rect 64259 200085 64287 200113
rect 64321 200085 64349 200113
rect 64383 200085 64411 200113
rect 64197 200023 64225 200051
rect 64259 200023 64287 200051
rect 64321 200023 64349 200051
rect 64383 200023 64411 200051
rect 64197 199961 64225 199989
rect 64259 199961 64287 199989
rect 64321 199961 64349 199989
rect 64383 199961 64411 199989
rect 64197 191147 64225 191175
rect 64259 191147 64287 191175
rect 64321 191147 64349 191175
rect 64383 191147 64411 191175
rect 64197 191085 64225 191113
rect 64259 191085 64287 191113
rect 64321 191085 64349 191113
rect 64383 191085 64411 191113
rect 64197 191023 64225 191051
rect 64259 191023 64287 191051
rect 64321 191023 64349 191051
rect 64383 191023 64411 191051
rect 64197 190961 64225 190989
rect 64259 190961 64287 190989
rect 64321 190961 64349 190989
rect 64383 190961 64411 190989
rect 64197 182147 64225 182175
rect 64259 182147 64287 182175
rect 64321 182147 64349 182175
rect 64383 182147 64411 182175
rect 64197 182085 64225 182113
rect 64259 182085 64287 182113
rect 64321 182085 64349 182113
rect 64383 182085 64411 182113
rect 64197 182023 64225 182051
rect 64259 182023 64287 182051
rect 64321 182023 64349 182051
rect 64383 182023 64411 182051
rect 64197 181961 64225 181989
rect 64259 181961 64287 181989
rect 64321 181961 64349 181989
rect 64383 181961 64411 181989
rect 64197 173147 64225 173175
rect 64259 173147 64287 173175
rect 64321 173147 64349 173175
rect 64383 173147 64411 173175
rect 64197 173085 64225 173113
rect 64259 173085 64287 173113
rect 64321 173085 64349 173113
rect 64383 173085 64411 173113
rect 64197 173023 64225 173051
rect 64259 173023 64287 173051
rect 64321 173023 64349 173051
rect 64383 173023 64411 173051
rect 64197 172961 64225 172989
rect 64259 172961 64287 172989
rect 64321 172961 64349 172989
rect 64383 172961 64411 172989
rect 64197 164147 64225 164175
rect 64259 164147 64287 164175
rect 64321 164147 64349 164175
rect 64383 164147 64411 164175
rect 64197 164085 64225 164113
rect 64259 164085 64287 164113
rect 64321 164085 64349 164113
rect 64383 164085 64411 164113
rect 64197 164023 64225 164051
rect 64259 164023 64287 164051
rect 64321 164023 64349 164051
rect 64383 164023 64411 164051
rect 64197 163961 64225 163989
rect 64259 163961 64287 163989
rect 64321 163961 64349 163989
rect 64383 163961 64411 163989
rect 64197 155147 64225 155175
rect 64259 155147 64287 155175
rect 64321 155147 64349 155175
rect 64383 155147 64411 155175
rect 64197 155085 64225 155113
rect 64259 155085 64287 155113
rect 64321 155085 64349 155113
rect 64383 155085 64411 155113
rect 64197 155023 64225 155051
rect 64259 155023 64287 155051
rect 64321 155023 64349 155051
rect 64383 155023 64411 155051
rect 64197 154961 64225 154989
rect 64259 154961 64287 154989
rect 64321 154961 64349 154989
rect 64383 154961 64411 154989
rect 64197 146147 64225 146175
rect 64259 146147 64287 146175
rect 64321 146147 64349 146175
rect 64383 146147 64411 146175
rect 64197 146085 64225 146113
rect 64259 146085 64287 146113
rect 64321 146085 64349 146113
rect 64383 146085 64411 146113
rect 64197 146023 64225 146051
rect 64259 146023 64287 146051
rect 64321 146023 64349 146051
rect 64383 146023 64411 146051
rect 64197 145961 64225 145989
rect 64259 145961 64287 145989
rect 64321 145961 64349 145989
rect 64383 145961 64411 145989
rect 64197 137147 64225 137175
rect 64259 137147 64287 137175
rect 64321 137147 64349 137175
rect 64383 137147 64411 137175
rect 64197 137085 64225 137113
rect 64259 137085 64287 137113
rect 64321 137085 64349 137113
rect 64383 137085 64411 137113
rect 64197 137023 64225 137051
rect 64259 137023 64287 137051
rect 64321 137023 64349 137051
rect 64383 137023 64411 137051
rect 64197 136961 64225 136989
rect 64259 136961 64287 136989
rect 64321 136961 64349 136989
rect 64383 136961 64411 136989
rect 64197 128147 64225 128175
rect 64259 128147 64287 128175
rect 64321 128147 64349 128175
rect 64383 128147 64411 128175
rect 64197 128085 64225 128113
rect 64259 128085 64287 128113
rect 64321 128085 64349 128113
rect 64383 128085 64411 128113
rect 64197 128023 64225 128051
rect 64259 128023 64287 128051
rect 64321 128023 64349 128051
rect 64383 128023 64411 128051
rect 64197 127961 64225 127989
rect 64259 127961 64287 127989
rect 64321 127961 64349 127989
rect 64383 127961 64411 127989
rect 64197 119147 64225 119175
rect 64259 119147 64287 119175
rect 64321 119147 64349 119175
rect 64383 119147 64411 119175
rect 64197 119085 64225 119113
rect 64259 119085 64287 119113
rect 64321 119085 64349 119113
rect 64383 119085 64411 119113
rect 64197 119023 64225 119051
rect 64259 119023 64287 119051
rect 64321 119023 64349 119051
rect 64383 119023 64411 119051
rect 64197 118961 64225 118989
rect 64259 118961 64287 118989
rect 64321 118961 64349 118989
rect 64383 118961 64411 118989
rect 64197 110147 64225 110175
rect 64259 110147 64287 110175
rect 64321 110147 64349 110175
rect 64383 110147 64411 110175
rect 64197 110085 64225 110113
rect 64259 110085 64287 110113
rect 64321 110085 64349 110113
rect 64383 110085 64411 110113
rect 64197 110023 64225 110051
rect 64259 110023 64287 110051
rect 64321 110023 64349 110051
rect 64383 110023 64411 110051
rect 64197 109961 64225 109989
rect 64259 109961 64287 109989
rect 64321 109961 64349 109989
rect 64383 109961 64411 109989
rect 64197 101147 64225 101175
rect 64259 101147 64287 101175
rect 64321 101147 64349 101175
rect 64383 101147 64411 101175
rect 64197 101085 64225 101113
rect 64259 101085 64287 101113
rect 64321 101085 64349 101113
rect 64383 101085 64411 101113
rect 64197 101023 64225 101051
rect 64259 101023 64287 101051
rect 64321 101023 64349 101051
rect 64383 101023 64411 101051
rect 64197 100961 64225 100989
rect 64259 100961 64287 100989
rect 64321 100961 64349 100989
rect 64383 100961 64411 100989
rect 64197 92147 64225 92175
rect 64259 92147 64287 92175
rect 64321 92147 64349 92175
rect 64383 92147 64411 92175
rect 64197 92085 64225 92113
rect 64259 92085 64287 92113
rect 64321 92085 64349 92113
rect 64383 92085 64411 92113
rect 64197 92023 64225 92051
rect 64259 92023 64287 92051
rect 64321 92023 64349 92051
rect 64383 92023 64411 92051
rect 64197 91961 64225 91989
rect 64259 91961 64287 91989
rect 64321 91961 64349 91989
rect 64383 91961 64411 91989
rect 64197 83147 64225 83175
rect 64259 83147 64287 83175
rect 64321 83147 64349 83175
rect 64383 83147 64411 83175
rect 64197 83085 64225 83113
rect 64259 83085 64287 83113
rect 64321 83085 64349 83113
rect 64383 83085 64411 83113
rect 64197 83023 64225 83051
rect 64259 83023 64287 83051
rect 64321 83023 64349 83051
rect 64383 83023 64411 83051
rect 64197 82961 64225 82989
rect 64259 82961 64287 82989
rect 64321 82961 64349 82989
rect 64383 82961 64411 82989
rect 64197 74147 64225 74175
rect 64259 74147 64287 74175
rect 64321 74147 64349 74175
rect 64383 74147 64411 74175
rect 64197 74085 64225 74113
rect 64259 74085 64287 74113
rect 64321 74085 64349 74113
rect 64383 74085 64411 74113
rect 64197 74023 64225 74051
rect 64259 74023 64287 74051
rect 64321 74023 64349 74051
rect 64383 74023 64411 74051
rect 64197 73961 64225 73989
rect 64259 73961 64287 73989
rect 64321 73961 64349 73989
rect 64383 73961 64411 73989
rect 64197 65147 64225 65175
rect 64259 65147 64287 65175
rect 64321 65147 64349 65175
rect 64383 65147 64411 65175
rect 64197 65085 64225 65113
rect 64259 65085 64287 65113
rect 64321 65085 64349 65113
rect 64383 65085 64411 65113
rect 64197 65023 64225 65051
rect 64259 65023 64287 65051
rect 64321 65023 64349 65051
rect 64383 65023 64411 65051
rect 64197 64961 64225 64989
rect 64259 64961 64287 64989
rect 64321 64961 64349 64989
rect 64383 64961 64411 64989
rect 64197 56147 64225 56175
rect 64259 56147 64287 56175
rect 64321 56147 64349 56175
rect 64383 56147 64411 56175
rect 64197 56085 64225 56113
rect 64259 56085 64287 56113
rect 64321 56085 64349 56113
rect 64383 56085 64411 56113
rect 64197 56023 64225 56051
rect 64259 56023 64287 56051
rect 64321 56023 64349 56051
rect 64383 56023 64411 56051
rect 64197 55961 64225 55989
rect 64259 55961 64287 55989
rect 64321 55961 64349 55989
rect 64383 55961 64411 55989
rect 64197 47147 64225 47175
rect 64259 47147 64287 47175
rect 64321 47147 64349 47175
rect 64383 47147 64411 47175
rect 64197 47085 64225 47113
rect 64259 47085 64287 47113
rect 64321 47085 64349 47113
rect 64383 47085 64411 47113
rect 64197 47023 64225 47051
rect 64259 47023 64287 47051
rect 64321 47023 64349 47051
rect 64383 47023 64411 47051
rect 64197 46961 64225 46989
rect 64259 46961 64287 46989
rect 64321 46961 64349 46989
rect 64383 46961 64411 46989
rect 64197 38147 64225 38175
rect 64259 38147 64287 38175
rect 64321 38147 64349 38175
rect 64383 38147 64411 38175
rect 64197 38085 64225 38113
rect 64259 38085 64287 38113
rect 64321 38085 64349 38113
rect 64383 38085 64411 38113
rect 64197 38023 64225 38051
rect 64259 38023 64287 38051
rect 64321 38023 64349 38051
rect 64383 38023 64411 38051
rect 64197 37961 64225 37989
rect 64259 37961 64287 37989
rect 64321 37961 64349 37989
rect 64383 37961 64411 37989
rect 64197 29147 64225 29175
rect 64259 29147 64287 29175
rect 64321 29147 64349 29175
rect 64383 29147 64411 29175
rect 64197 29085 64225 29113
rect 64259 29085 64287 29113
rect 64321 29085 64349 29113
rect 64383 29085 64411 29113
rect 64197 29023 64225 29051
rect 64259 29023 64287 29051
rect 64321 29023 64349 29051
rect 64383 29023 64411 29051
rect 64197 28961 64225 28989
rect 64259 28961 64287 28989
rect 64321 28961 64349 28989
rect 64383 28961 64411 28989
rect 64197 20147 64225 20175
rect 64259 20147 64287 20175
rect 64321 20147 64349 20175
rect 64383 20147 64411 20175
rect 64197 20085 64225 20113
rect 64259 20085 64287 20113
rect 64321 20085 64349 20113
rect 64383 20085 64411 20113
rect 64197 20023 64225 20051
rect 64259 20023 64287 20051
rect 64321 20023 64349 20051
rect 64383 20023 64411 20051
rect 64197 19961 64225 19989
rect 64259 19961 64287 19989
rect 64321 19961 64349 19989
rect 64383 19961 64411 19989
rect 64197 11147 64225 11175
rect 64259 11147 64287 11175
rect 64321 11147 64349 11175
rect 64383 11147 64411 11175
rect 64197 11085 64225 11113
rect 64259 11085 64287 11113
rect 64321 11085 64349 11113
rect 64383 11085 64411 11113
rect 64197 11023 64225 11051
rect 64259 11023 64287 11051
rect 64321 11023 64349 11051
rect 64383 11023 64411 11051
rect 64197 10961 64225 10989
rect 64259 10961 64287 10989
rect 64321 10961 64349 10989
rect 64383 10961 64411 10989
rect 64197 2147 64225 2175
rect 64259 2147 64287 2175
rect 64321 2147 64349 2175
rect 64383 2147 64411 2175
rect 64197 2085 64225 2113
rect 64259 2085 64287 2113
rect 64321 2085 64349 2113
rect 64383 2085 64411 2113
rect 64197 2023 64225 2051
rect 64259 2023 64287 2051
rect 64321 2023 64349 2051
rect 64383 2023 64411 2051
rect 64197 1961 64225 1989
rect 64259 1961 64287 1989
rect 64321 1961 64349 1989
rect 64383 1961 64411 1989
rect 64197 -108 64225 -80
rect 64259 -108 64287 -80
rect 64321 -108 64349 -80
rect 64383 -108 64411 -80
rect 64197 -170 64225 -142
rect 64259 -170 64287 -142
rect 64321 -170 64349 -142
rect 64383 -170 64411 -142
rect 64197 -232 64225 -204
rect 64259 -232 64287 -204
rect 64321 -232 64349 -204
rect 64383 -232 64411 -204
rect 64197 -294 64225 -266
rect 64259 -294 64287 -266
rect 64321 -294 64349 -266
rect 64383 -294 64411 -266
rect 66057 299058 66085 299086
rect 66119 299058 66147 299086
rect 66181 299058 66209 299086
rect 66243 299058 66271 299086
rect 66057 298996 66085 299024
rect 66119 298996 66147 299024
rect 66181 298996 66209 299024
rect 66243 298996 66271 299024
rect 66057 298934 66085 298962
rect 66119 298934 66147 298962
rect 66181 298934 66209 298962
rect 66243 298934 66271 298962
rect 66057 298872 66085 298900
rect 66119 298872 66147 298900
rect 66181 298872 66209 298900
rect 66243 298872 66271 298900
rect 66057 293147 66085 293175
rect 66119 293147 66147 293175
rect 66181 293147 66209 293175
rect 66243 293147 66271 293175
rect 66057 293085 66085 293113
rect 66119 293085 66147 293113
rect 66181 293085 66209 293113
rect 66243 293085 66271 293113
rect 66057 293023 66085 293051
rect 66119 293023 66147 293051
rect 66181 293023 66209 293051
rect 66243 293023 66271 293051
rect 66057 292961 66085 292989
rect 66119 292961 66147 292989
rect 66181 292961 66209 292989
rect 66243 292961 66271 292989
rect 66057 284147 66085 284175
rect 66119 284147 66147 284175
rect 66181 284147 66209 284175
rect 66243 284147 66271 284175
rect 66057 284085 66085 284113
rect 66119 284085 66147 284113
rect 66181 284085 66209 284113
rect 66243 284085 66271 284113
rect 66057 284023 66085 284051
rect 66119 284023 66147 284051
rect 66181 284023 66209 284051
rect 66243 284023 66271 284051
rect 66057 283961 66085 283989
rect 66119 283961 66147 283989
rect 66181 283961 66209 283989
rect 66243 283961 66271 283989
rect 66057 275147 66085 275175
rect 66119 275147 66147 275175
rect 66181 275147 66209 275175
rect 66243 275147 66271 275175
rect 66057 275085 66085 275113
rect 66119 275085 66147 275113
rect 66181 275085 66209 275113
rect 66243 275085 66271 275113
rect 66057 275023 66085 275051
rect 66119 275023 66147 275051
rect 66181 275023 66209 275051
rect 66243 275023 66271 275051
rect 66057 274961 66085 274989
rect 66119 274961 66147 274989
rect 66181 274961 66209 274989
rect 66243 274961 66271 274989
rect 66057 266147 66085 266175
rect 66119 266147 66147 266175
rect 66181 266147 66209 266175
rect 66243 266147 66271 266175
rect 66057 266085 66085 266113
rect 66119 266085 66147 266113
rect 66181 266085 66209 266113
rect 66243 266085 66271 266113
rect 66057 266023 66085 266051
rect 66119 266023 66147 266051
rect 66181 266023 66209 266051
rect 66243 266023 66271 266051
rect 66057 265961 66085 265989
rect 66119 265961 66147 265989
rect 66181 265961 66209 265989
rect 66243 265961 66271 265989
rect 66057 257147 66085 257175
rect 66119 257147 66147 257175
rect 66181 257147 66209 257175
rect 66243 257147 66271 257175
rect 66057 257085 66085 257113
rect 66119 257085 66147 257113
rect 66181 257085 66209 257113
rect 66243 257085 66271 257113
rect 66057 257023 66085 257051
rect 66119 257023 66147 257051
rect 66181 257023 66209 257051
rect 66243 257023 66271 257051
rect 66057 256961 66085 256989
rect 66119 256961 66147 256989
rect 66181 256961 66209 256989
rect 66243 256961 66271 256989
rect 66057 248147 66085 248175
rect 66119 248147 66147 248175
rect 66181 248147 66209 248175
rect 66243 248147 66271 248175
rect 66057 248085 66085 248113
rect 66119 248085 66147 248113
rect 66181 248085 66209 248113
rect 66243 248085 66271 248113
rect 66057 248023 66085 248051
rect 66119 248023 66147 248051
rect 66181 248023 66209 248051
rect 66243 248023 66271 248051
rect 66057 247961 66085 247989
rect 66119 247961 66147 247989
rect 66181 247961 66209 247989
rect 66243 247961 66271 247989
rect 66057 239147 66085 239175
rect 66119 239147 66147 239175
rect 66181 239147 66209 239175
rect 66243 239147 66271 239175
rect 66057 239085 66085 239113
rect 66119 239085 66147 239113
rect 66181 239085 66209 239113
rect 66243 239085 66271 239113
rect 66057 239023 66085 239051
rect 66119 239023 66147 239051
rect 66181 239023 66209 239051
rect 66243 239023 66271 239051
rect 66057 238961 66085 238989
rect 66119 238961 66147 238989
rect 66181 238961 66209 238989
rect 66243 238961 66271 238989
rect 66057 230147 66085 230175
rect 66119 230147 66147 230175
rect 66181 230147 66209 230175
rect 66243 230147 66271 230175
rect 66057 230085 66085 230113
rect 66119 230085 66147 230113
rect 66181 230085 66209 230113
rect 66243 230085 66271 230113
rect 66057 230023 66085 230051
rect 66119 230023 66147 230051
rect 66181 230023 66209 230051
rect 66243 230023 66271 230051
rect 66057 229961 66085 229989
rect 66119 229961 66147 229989
rect 66181 229961 66209 229989
rect 66243 229961 66271 229989
rect 66057 221147 66085 221175
rect 66119 221147 66147 221175
rect 66181 221147 66209 221175
rect 66243 221147 66271 221175
rect 66057 221085 66085 221113
rect 66119 221085 66147 221113
rect 66181 221085 66209 221113
rect 66243 221085 66271 221113
rect 66057 221023 66085 221051
rect 66119 221023 66147 221051
rect 66181 221023 66209 221051
rect 66243 221023 66271 221051
rect 66057 220961 66085 220989
rect 66119 220961 66147 220989
rect 66181 220961 66209 220989
rect 66243 220961 66271 220989
rect 66057 212147 66085 212175
rect 66119 212147 66147 212175
rect 66181 212147 66209 212175
rect 66243 212147 66271 212175
rect 66057 212085 66085 212113
rect 66119 212085 66147 212113
rect 66181 212085 66209 212113
rect 66243 212085 66271 212113
rect 66057 212023 66085 212051
rect 66119 212023 66147 212051
rect 66181 212023 66209 212051
rect 66243 212023 66271 212051
rect 66057 211961 66085 211989
rect 66119 211961 66147 211989
rect 66181 211961 66209 211989
rect 66243 211961 66271 211989
rect 66057 203147 66085 203175
rect 66119 203147 66147 203175
rect 66181 203147 66209 203175
rect 66243 203147 66271 203175
rect 66057 203085 66085 203113
rect 66119 203085 66147 203113
rect 66181 203085 66209 203113
rect 66243 203085 66271 203113
rect 66057 203023 66085 203051
rect 66119 203023 66147 203051
rect 66181 203023 66209 203051
rect 66243 203023 66271 203051
rect 66057 202961 66085 202989
rect 66119 202961 66147 202989
rect 66181 202961 66209 202989
rect 66243 202961 66271 202989
rect 66057 194147 66085 194175
rect 66119 194147 66147 194175
rect 66181 194147 66209 194175
rect 66243 194147 66271 194175
rect 66057 194085 66085 194113
rect 66119 194085 66147 194113
rect 66181 194085 66209 194113
rect 66243 194085 66271 194113
rect 66057 194023 66085 194051
rect 66119 194023 66147 194051
rect 66181 194023 66209 194051
rect 66243 194023 66271 194051
rect 66057 193961 66085 193989
rect 66119 193961 66147 193989
rect 66181 193961 66209 193989
rect 66243 193961 66271 193989
rect 66057 185147 66085 185175
rect 66119 185147 66147 185175
rect 66181 185147 66209 185175
rect 66243 185147 66271 185175
rect 66057 185085 66085 185113
rect 66119 185085 66147 185113
rect 66181 185085 66209 185113
rect 66243 185085 66271 185113
rect 66057 185023 66085 185051
rect 66119 185023 66147 185051
rect 66181 185023 66209 185051
rect 66243 185023 66271 185051
rect 66057 184961 66085 184989
rect 66119 184961 66147 184989
rect 66181 184961 66209 184989
rect 66243 184961 66271 184989
rect 66057 176147 66085 176175
rect 66119 176147 66147 176175
rect 66181 176147 66209 176175
rect 66243 176147 66271 176175
rect 66057 176085 66085 176113
rect 66119 176085 66147 176113
rect 66181 176085 66209 176113
rect 66243 176085 66271 176113
rect 66057 176023 66085 176051
rect 66119 176023 66147 176051
rect 66181 176023 66209 176051
rect 66243 176023 66271 176051
rect 66057 175961 66085 175989
rect 66119 175961 66147 175989
rect 66181 175961 66209 175989
rect 66243 175961 66271 175989
rect 66057 167147 66085 167175
rect 66119 167147 66147 167175
rect 66181 167147 66209 167175
rect 66243 167147 66271 167175
rect 66057 167085 66085 167113
rect 66119 167085 66147 167113
rect 66181 167085 66209 167113
rect 66243 167085 66271 167113
rect 66057 167023 66085 167051
rect 66119 167023 66147 167051
rect 66181 167023 66209 167051
rect 66243 167023 66271 167051
rect 66057 166961 66085 166989
rect 66119 166961 66147 166989
rect 66181 166961 66209 166989
rect 66243 166961 66271 166989
rect 66057 158147 66085 158175
rect 66119 158147 66147 158175
rect 66181 158147 66209 158175
rect 66243 158147 66271 158175
rect 66057 158085 66085 158113
rect 66119 158085 66147 158113
rect 66181 158085 66209 158113
rect 66243 158085 66271 158113
rect 66057 158023 66085 158051
rect 66119 158023 66147 158051
rect 66181 158023 66209 158051
rect 66243 158023 66271 158051
rect 66057 157961 66085 157989
rect 66119 157961 66147 157989
rect 66181 157961 66209 157989
rect 66243 157961 66271 157989
rect 66057 149147 66085 149175
rect 66119 149147 66147 149175
rect 66181 149147 66209 149175
rect 66243 149147 66271 149175
rect 66057 149085 66085 149113
rect 66119 149085 66147 149113
rect 66181 149085 66209 149113
rect 66243 149085 66271 149113
rect 66057 149023 66085 149051
rect 66119 149023 66147 149051
rect 66181 149023 66209 149051
rect 66243 149023 66271 149051
rect 66057 148961 66085 148989
rect 66119 148961 66147 148989
rect 66181 148961 66209 148989
rect 66243 148961 66271 148989
rect 66057 140147 66085 140175
rect 66119 140147 66147 140175
rect 66181 140147 66209 140175
rect 66243 140147 66271 140175
rect 66057 140085 66085 140113
rect 66119 140085 66147 140113
rect 66181 140085 66209 140113
rect 66243 140085 66271 140113
rect 66057 140023 66085 140051
rect 66119 140023 66147 140051
rect 66181 140023 66209 140051
rect 66243 140023 66271 140051
rect 66057 139961 66085 139989
rect 66119 139961 66147 139989
rect 66181 139961 66209 139989
rect 66243 139961 66271 139989
rect 66057 131147 66085 131175
rect 66119 131147 66147 131175
rect 66181 131147 66209 131175
rect 66243 131147 66271 131175
rect 66057 131085 66085 131113
rect 66119 131085 66147 131113
rect 66181 131085 66209 131113
rect 66243 131085 66271 131113
rect 66057 131023 66085 131051
rect 66119 131023 66147 131051
rect 66181 131023 66209 131051
rect 66243 131023 66271 131051
rect 66057 130961 66085 130989
rect 66119 130961 66147 130989
rect 66181 130961 66209 130989
rect 66243 130961 66271 130989
rect 66057 122147 66085 122175
rect 66119 122147 66147 122175
rect 66181 122147 66209 122175
rect 66243 122147 66271 122175
rect 66057 122085 66085 122113
rect 66119 122085 66147 122113
rect 66181 122085 66209 122113
rect 66243 122085 66271 122113
rect 66057 122023 66085 122051
rect 66119 122023 66147 122051
rect 66181 122023 66209 122051
rect 66243 122023 66271 122051
rect 66057 121961 66085 121989
rect 66119 121961 66147 121989
rect 66181 121961 66209 121989
rect 66243 121961 66271 121989
rect 66057 113147 66085 113175
rect 66119 113147 66147 113175
rect 66181 113147 66209 113175
rect 66243 113147 66271 113175
rect 66057 113085 66085 113113
rect 66119 113085 66147 113113
rect 66181 113085 66209 113113
rect 66243 113085 66271 113113
rect 66057 113023 66085 113051
rect 66119 113023 66147 113051
rect 66181 113023 66209 113051
rect 66243 113023 66271 113051
rect 66057 112961 66085 112989
rect 66119 112961 66147 112989
rect 66181 112961 66209 112989
rect 66243 112961 66271 112989
rect 66057 104147 66085 104175
rect 66119 104147 66147 104175
rect 66181 104147 66209 104175
rect 66243 104147 66271 104175
rect 66057 104085 66085 104113
rect 66119 104085 66147 104113
rect 66181 104085 66209 104113
rect 66243 104085 66271 104113
rect 66057 104023 66085 104051
rect 66119 104023 66147 104051
rect 66181 104023 66209 104051
rect 66243 104023 66271 104051
rect 66057 103961 66085 103989
rect 66119 103961 66147 103989
rect 66181 103961 66209 103989
rect 66243 103961 66271 103989
rect 66057 95147 66085 95175
rect 66119 95147 66147 95175
rect 66181 95147 66209 95175
rect 66243 95147 66271 95175
rect 66057 95085 66085 95113
rect 66119 95085 66147 95113
rect 66181 95085 66209 95113
rect 66243 95085 66271 95113
rect 66057 95023 66085 95051
rect 66119 95023 66147 95051
rect 66181 95023 66209 95051
rect 66243 95023 66271 95051
rect 66057 94961 66085 94989
rect 66119 94961 66147 94989
rect 66181 94961 66209 94989
rect 66243 94961 66271 94989
rect 66057 86147 66085 86175
rect 66119 86147 66147 86175
rect 66181 86147 66209 86175
rect 66243 86147 66271 86175
rect 66057 86085 66085 86113
rect 66119 86085 66147 86113
rect 66181 86085 66209 86113
rect 66243 86085 66271 86113
rect 66057 86023 66085 86051
rect 66119 86023 66147 86051
rect 66181 86023 66209 86051
rect 66243 86023 66271 86051
rect 66057 85961 66085 85989
rect 66119 85961 66147 85989
rect 66181 85961 66209 85989
rect 66243 85961 66271 85989
rect 66057 77147 66085 77175
rect 66119 77147 66147 77175
rect 66181 77147 66209 77175
rect 66243 77147 66271 77175
rect 66057 77085 66085 77113
rect 66119 77085 66147 77113
rect 66181 77085 66209 77113
rect 66243 77085 66271 77113
rect 66057 77023 66085 77051
rect 66119 77023 66147 77051
rect 66181 77023 66209 77051
rect 66243 77023 66271 77051
rect 66057 76961 66085 76989
rect 66119 76961 66147 76989
rect 66181 76961 66209 76989
rect 66243 76961 66271 76989
rect 66057 68147 66085 68175
rect 66119 68147 66147 68175
rect 66181 68147 66209 68175
rect 66243 68147 66271 68175
rect 66057 68085 66085 68113
rect 66119 68085 66147 68113
rect 66181 68085 66209 68113
rect 66243 68085 66271 68113
rect 66057 68023 66085 68051
rect 66119 68023 66147 68051
rect 66181 68023 66209 68051
rect 66243 68023 66271 68051
rect 66057 67961 66085 67989
rect 66119 67961 66147 67989
rect 66181 67961 66209 67989
rect 66243 67961 66271 67989
rect 66057 59147 66085 59175
rect 66119 59147 66147 59175
rect 66181 59147 66209 59175
rect 66243 59147 66271 59175
rect 66057 59085 66085 59113
rect 66119 59085 66147 59113
rect 66181 59085 66209 59113
rect 66243 59085 66271 59113
rect 66057 59023 66085 59051
rect 66119 59023 66147 59051
rect 66181 59023 66209 59051
rect 66243 59023 66271 59051
rect 66057 58961 66085 58989
rect 66119 58961 66147 58989
rect 66181 58961 66209 58989
rect 66243 58961 66271 58989
rect 66057 50147 66085 50175
rect 66119 50147 66147 50175
rect 66181 50147 66209 50175
rect 66243 50147 66271 50175
rect 66057 50085 66085 50113
rect 66119 50085 66147 50113
rect 66181 50085 66209 50113
rect 66243 50085 66271 50113
rect 66057 50023 66085 50051
rect 66119 50023 66147 50051
rect 66181 50023 66209 50051
rect 66243 50023 66271 50051
rect 66057 49961 66085 49989
rect 66119 49961 66147 49989
rect 66181 49961 66209 49989
rect 66243 49961 66271 49989
rect 66057 41147 66085 41175
rect 66119 41147 66147 41175
rect 66181 41147 66209 41175
rect 66243 41147 66271 41175
rect 66057 41085 66085 41113
rect 66119 41085 66147 41113
rect 66181 41085 66209 41113
rect 66243 41085 66271 41113
rect 66057 41023 66085 41051
rect 66119 41023 66147 41051
rect 66181 41023 66209 41051
rect 66243 41023 66271 41051
rect 66057 40961 66085 40989
rect 66119 40961 66147 40989
rect 66181 40961 66209 40989
rect 66243 40961 66271 40989
rect 66057 32147 66085 32175
rect 66119 32147 66147 32175
rect 66181 32147 66209 32175
rect 66243 32147 66271 32175
rect 66057 32085 66085 32113
rect 66119 32085 66147 32113
rect 66181 32085 66209 32113
rect 66243 32085 66271 32113
rect 66057 32023 66085 32051
rect 66119 32023 66147 32051
rect 66181 32023 66209 32051
rect 66243 32023 66271 32051
rect 66057 31961 66085 31989
rect 66119 31961 66147 31989
rect 66181 31961 66209 31989
rect 66243 31961 66271 31989
rect 66057 23147 66085 23175
rect 66119 23147 66147 23175
rect 66181 23147 66209 23175
rect 66243 23147 66271 23175
rect 66057 23085 66085 23113
rect 66119 23085 66147 23113
rect 66181 23085 66209 23113
rect 66243 23085 66271 23113
rect 66057 23023 66085 23051
rect 66119 23023 66147 23051
rect 66181 23023 66209 23051
rect 66243 23023 66271 23051
rect 66057 22961 66085 22989
rect 66119 22961 66147 22989
rect 66181 22961 66209 22989
rect 66243 22961 66271 22989
rect 66057 14147 66085 14175
rect 66119 14147 66147 14175
rect 66181 14147 66209 14175
rect 66243 14147 66271 14175
rect 66057 14085 66085 14113
rect 66119 14085 66147 14113
rect 66181 14085 66209 14113
rect 66243 14085 66271 14113
rect 66057 14023 66085 14051
rect 66119 14023 66147 14051
rect 66181 14023 66209 14051
rect 66243 14023 66271 14051
rect 66057 13961 66085 13989
rect 66119 13961 66147 13989
rect 66181 13961 66209 13989
rect 66243 13961 66271 13989
rect 66057 5147 66085 5175
rect 66119 5147 66147 5175
rect 66181 5147 66209 5175
rect 66243 5147 66271 5175
rect 66057 5085 66085 5113
rect 66119 5085 66147 5113
rect 66181 5085 66209 5113
rect 66243 5085 66271 5113
rect 66057 5023 66085 5051
rect 66119 5023 66147 5051
rect 66181 5023 66209 5051
rect 66243 5023 66271 5051
rect 66057 4961 66085 4989
rect 66119 4961 66147 4989
rect 66181 4961 66209 4989
rect 66243 4961 66271 4989
rect 66057 -588 66085 -560
rect 66119 -588 66147 -560
rect 66181 -588 66209 -560
rect 66243 -588 66271 -560
rect 66057 -650 66085 -622
rect 66119 -650 66147 -622
rect 66181 -650 66209 -622
rect 66243 -650 66271 -622
rect 66057 -712 66085 -684
rect 66119 -712 66147 -684
rect 66181 -712 66209 -684
rect 66243 -712 66271 -684
rect 66057 -774 66085 -746
rect 66119 -774 66147 -746
rect 66181 -774 66209 -746
rect 66243 -774 66271 -746
rect 79557 298578 79585 298606
rect 79619 298578 79647 298606
rect 79681 298578 79709 298606
rect 79743 298578 79771 298606
rect 79557 298516 79585 298544
rect 79619 298516 79647 298544
rect 79681 298516 79709 298544
rect 79743 298516 79771 298544
rect 79557 298454 79585 298482
rect 79619 298454 79647 298482
rect 79681 298454 79709 298482
rect 79743 298454 79771 298482
rect 79557 298392 79585 298420
rect 79619 298392 79647 298420
rect 79681 298392 79709 298420
rect 79743 298392 79771 298420
rect 79557 290147 79585 290175
rect 79619 290147 79647 290175
rect 79681 290147 79709 290175
rect 79743 290147 79771 290175
rect 79557 290085 79585 290113
rect 79619 290085 79647 290113
rect 79681 290085 79709 290113
rect 79743 290085 79771 290113
rect 79557 290023 79585 290051
rect 79619 290023 79647 290051
rect 79681 290023 79709 290051
rect 79743 290023 79771 290051
rect 79557 289961 79585 289989
rect 79619 289961 79647 289989
rect 79681 289961 79709 289989
rect 79743 289961 79771 289989
rect 79557 281147 79585 281175
rect 79619 281147 79647 281175
rect 79681 281147 79709 281175
rect 79743 281147 79771 281175
rect 79557 281085 79585 281113
rect 79619 281085 79647 281113
rect 79681 281085 79709 281113
rect 79743 281085 79771 281113
rect 79557 281023 79585 281051
rect 79619 281023 79647 281051
rect 79681 281023 79709 281051
rect 79743 281023 79771 281051
rect 79557 280961 79585 280989
rect 79619 280961 79647 280989
rect 79681 280961 79709 280989
rect 79743 280961 79771 280989
rect 79557 272147 79585 272175
rect 79619 272147 79647 272175
rect 79681 272147 79709 272175
rect 79743 272147 79771 272175
rect 79557 272085 79585 272113
rect 79619 272085 79647 272113
rect 79681 272085 79709 272113
rect 79743 272085 79771 272113
rect 79557 272023 79585 272051
rect 79619 272023 79647 272051
rect 79681 272023 79709 272051
rect 79743 272023 79771 272051
rect 79557 271961 79585 271989
rect 79619 271961 79647 271989
rect 79681 271961 79709 271989
rect 79743 271961 79771 271989
rect 79557 263147 79585 263175
rect 79619 263147 79647 263175
rect 79681 263147 79709 263175
rect 79743 263147 79771 263175
rect 79557 263085 79585 263113
rect 79619 263085 79647 263113
rect 79681 263085 79709 263113
rect 79743 263085 79771 263113
rect 79557 263023 79585 263051
rect 79619 263023 79647 263051
rect 79681 263023 79709 263051
rect 79743 263023 79771 263051
rect 79557 262961 79585 262989
rect 79619 262961 79647 262989
rect 79681 262961 79709 262989
rect 79743 262961 79771 262989
rect 79557 254147 79585 254175
rect 79619 254147 79647 254175
rect 79681 254147 79709 254175
rect 79743 254147 79771 254175
rect 79557 254085 79585 254113
rect 79619 254085 79647 254113
rect 79681 254085 79709 254113
rect 79743 254085 79771 254113
rect 79557 254023 79585 254051
rect 79619 254023 79647 254051
rect 79681 254023 79709 254051
rect 79743 254023 79771 254051
rect 79557 253961 79585 253989
rect 79619 253961 79647 253989
rect 79681 253961 79709 253989
rect 79743 253961 79771 253989
rect 79557 245147 79585 245175
rect 79619 245147 79647 245175
rect 79681 245147 79709 245175
rect 79743 245147 79771 245175
rect 79557 245085 79585 245113
rect 79619 245085 79647 245113
rect 79681 245085 79709 245113
rect 79743 245085 79771 245113
rect 79557 245023 79585 245051
rect 79619 245023 79647 245051
rect 79681 245023 79709 245051
rect 79743 245023 79771 245051
rect 79557 244961 79585 244989
rect 79619 244961 79647 244989
rect 79681 244961 79709 244989
rect 79743 244961 79771 244989
rect 79557 236147 79585 236175
rect 79619 236147 79647 236175
rect 79681 236147 79709 236175
rect 79743 236147 79771 236175
rect 79557 236085 79585 236113
rect 79619 236085 79647 236113
rect 79681 236085 79709 236113
rect 79743 236085 79771 236113
rect 79557 236023 79585 236051
rect 79619 236023 79647 236051
rect 79681 236023 79709 236051
rect 79743 236023 79771 236051
rect 79557 235961 79585 235989
rect 79619 235961 79647 235989
rect 79681 235961 79709 235989
rect 79743 235961 79771 235989
rect 79557 227147 79585 227175
rect 79619 227147 79647 227175
rect 79681 227147 79709 227175
rect 79743 227147 79771 227175
rect 79557 227085 79585 227113
rect 79619 227085 79647 227113
rect 79681 227085 79709 227113
rect 79743 227085 79771 227113
rect 79557 227023 79585 227051
rect 79619 227023 79647 227051
rect 79681 227023 79709 227051
rect 79743 227023 79771 227051
rect 79557 226961 79585 226989
rect 79619 226961 79647 226989
rect 79681 226961 79709 226989
rect 79743 226961 79771 226989
rect 79557 218147 79585 218175
rect 79619 218147 79647 218175
rect 79681 218147 79709 218175
rect 79743 218147 79771 218175
rect 79557 218085 79585 218113
rect 79619 218085 79647 218113
rect 79681 218085 79709 218113
rect 79743 218085 79771 218113
rect 79557 218023 79585 218051
rect 79619 218023 79647 218051
rect 79681 218023 79709 218051
rect 79743 218023 79771 218051
rect 79557 217961 79585 217989
rect 79619 217961 79647 217989
rect 79681 217961 79709 217989
rect 79743 217961 79771 217989
rect 79557 209147 79585 209175
rect 79619 209147 79647 209175
rect 79681 209147 79709 209175
rect 79743 209147 79771 209175
rect 79557 209085 79585 209113
rect 79619 209085 79647 209113
rect 79681 209085 79709 209113
rect 79743 209085 79771 209113
rect 79557 209023 79585 209051
rect 79619 209023 79647 209051
rect 79681 209023 79709 209051
rect 79743 209023 79771 209051
rect 79557 208961 79585 208989
rect 79619 208961 79647 208989
rect 79681 208961 79709 208989
rect 79743 208961 79771 208989
rect 79557 200147 79585 200175
rect 79619 200147 79647 200175
rect 79681 200147 79709 200175
rect 79743 200147 79771 200175
rect 79557 200085 79585 200113
rect 79619 200085 79647 200113
rect 79681 200085 79709 200113
rect 79743 200085 79771 200113
rect 79557 200023 79585 200051
rect 79619 200023 79647 200051
rect 79681 200023 79709 200051
rect 79743 200023 79771 200051
rect 79557 199961 79585 199989
rect 79619 199961 79647 199989
rect 79681 199961 79709 199989
rect 79743 199961 79771 199989
rect 79557 191147 79585 191175
rect 79619 191147 79647 191175
rect 79681 191147 79709 191175
rect 79743 191147 79771 191175
rect 79557 191085 79585 191113
rect 79619 191085 79647 191113
rect 79681 191085 79709 191113
rect 79743 191085 79771 191113
rect 79557 191023 79585 191051
rect 79619 191023 79647 191051
rect 79681 191023 79709 191051
rect 79743 191023 79771 191051
rect 79557 190961 79585 190989
rect 79619 190961 79647 190989
rect 79681 190961 79709 190989
rect 79743 190961 79771 190989
rect 79557 182147 79585 182175
rect 79619 182147 79647 182175
rect 79681 182147 79709 182175
rect 79743 182147 79771 182175
rect 79557 182085 79585 182113
rect 79619 182085 79647 182113
rect 79681 182085 79709 182113
rect 79743 182085 79771 182113
rect 79557 182023 79585 182051
rect 79619 182023 79647 182051
rect 79681 182023 79709 182051
rect 79743 182023 79771 182051
rect 79557 181961 79585 181989
rect 79619 181961 79647 181989
rect 79681 181961 79709 181989
rect 79743 181961 79771 181989
rect 79557 173147 79585 173175
rect 79619 173147 79647 173175
rect 79681 173147 79709 173175
rect 79743 173147 79771 173175
rect 79557 173085 79585 173113
rect 79619 173085 79647 173113
rect 79681 173085 79709 173113
rect 79743 173085 79771 173113
rect 79557 173023 79585 173051
rect 79619 173023 79647 173051
rect 79681 173023 79709 173051
rect 79743 173023 79771 173051
rect 79557 172961 79585 172989
rect 79619 172961 79647 172989
rect 79681 172961 79709 172989
rect 79743 172961 79771 172989
rect 79557 164147 79585 164175
rect 79619 164147 79647 164175
rect 79681 164147 79709 164175
rect 79743 164147 79771 164175
rect 79557 164085 79585 164113
rect 79619 164085 79647 164113
rect 79681 164085 79709 164113
rect 79743 164085 79771 164113
rect 79557 164023 79585 164051
rect 79619 164023 79647 164051
rect 79681 164023 79709 164051
rect 79743 164023 79771 164051
rect 79557 163961 79585 163989
rect 79619 163961 79647 163989
rect 79681 163961 79709 163989
rect 79743 163961 79771 163989
rect 79557 155147 79585 155175
rect 79619 155147 79647 155175
rect 79681 155147 79709 155175
rect 79743 155147 79771 155175
rect 79557 155085 79585 155113
rect 79619 155085 79647 155113
rect 79681 155085 79709 155113
rect 79743 155085 79771 155113
rect 79557 155023 79585 155051
rect 79619 155023 79647 155051
rect 79681 155023 79709 155051
rect 79743 155023 79771 155051
rect 79557 154961 79585 154989
rect 79619 154961 79647 154989
rect 79681 154961 79709 154989
rect 79743 154961 79771 154989
rect 79557 146147 79585 146175
rect 79619 146147 79647 146175
rect 79681 146147 79709 146175
rect 79743 146147 79771 146175
rect 79557 146085 79585 146113
rect 79619 146085 79647 146113
rect 79681 146085 79709 146113
rect 79743 146085 79771 146113
rect 79557 146023 79585 146051
rect 79619 146023 79647 146051
rect 79681 146023 79709 146051
rect 79743 146023 79771 146051
rect 79557 145961 79585 145989
rect 79619 145961 79647 145989
rect 79681 145961 79709 145989
rect 79743 145961 79771 145989
rect 79557 137147 79585 137175
rect 79619 137147 79647 137175
rect 79681 137147 79709 137175
rect 79743 137147 79771 137175
rect 79557 137085 79585 137113
rect 79619 137085 79647 137113
rect 79681 137085 79709 137113
rect 79743 137085 79771 137113
rect 79557 137023 79585 137051
rect 79619 137023 79647 137051
rect 79681 137023 79709 137051
rect 79743 137023 79771 137051
rect 79557 136961 79585 136989
rect 79619 136961 79647 136989
rect 79681 136961 79709 136989
rect 79743 136961 79771 136989
rect 79557 128147 79585 128175
rect 79619 128147 79647 128175
rect 79681 128147 79709 128175
rect 79743 128147 79771 128175
rect 79557 128085 79585 128113
rect 79619 128085 79647 128113
rect 79681 128085 79709 128113
rect 79743 128085 79771 128113
rect 79557 128023 79585 128051
rect 79619 128023 79647 128051
rect 79681 128023 79709 128051
rect 79743 128023 79771 128051
rect 79557 127961 79585 127989
rect 79619 127961 79647 127989
rect 79681 127961 79709 127989
rect 79743 127961 79771 127989
rect 79557 119147 79585 119175
rect 79619 119147 79647 119175
rect 79681 119147 79709 119175
rect 79743 119147 79771 119175
rect 79557 119085 79585 119113
rect 79619 119085 79647 119113
rect 79681 119085 79709 119113
rect 79743 119085 79771 119113
rect 79557 119023 79585 119051
rect 79619 119023 79647 119051
rect 79681 119023 79709 119051
rect 79743 119023 79771 119051
rect 79557 118961 79585 118989
rect 79619 118961 79647 118989
rect 79681 118961 79709 118989
rect 79743 118961 79771 118989
rect 79557 110147 79585 110175
rect 79619 110147 79647 110175
rect 79681 110147 79709 110175
rect 79743 110147 79771 110175
rect 79557 110085 79585 110113
rect 79619 110085 79647 110113
rect 79681 110085 79709 110113
rect 79743 110085 79771 110113
rect 79557 110023 79585 110051
rect 79619 110023 79647 110051
rect 79681 110023 79709 110051
rect 79743 110023 79771 110051
rect 79557 109961 79585 109989
rect 79619 109961 79647 109989
rect 79681 109961 79709 109989
rect 79743 109961 79771 109989
rect 79557 101147 79585 101175
rect 79619 101147 79647 101175
rect 79681 101147 79709 101175
rect 79743 101147 79771 101175
rect 79557 101085 79585 101113
rect 79619 101085 79647 101113
rect 79681 101085 79709 101113
rect 79743 101085 79771 101113
rect 79557 101023 79585 101051
rect 79619 101023 79647 101051
rect 79681 101023 79709 101051
rect 79743 101023 79771 101051
rect 79557 100961 79585 100989
rect 79619 100961 79647 100989
rect 79681 100961 79709 100989
rect 79743 100961 79771 100989
rect 79557 92147 79585 92175
rect 79619 92147 79647 92175
rect 79681 92147 79709 92175
rect 79743 92147 79771 92175
rect 79557 92085 79585 92113
rect 79619 92085 79647 92113
rect 79681 92085 79709 92113
rect 79743 92085 79771 92113
rect 79557 92023 79585 92051
rect 79619 92023 79647 92051
rect 79681 92023 79709 92051
rect 79743 92023 79771 92051
rect 79557 91961 79585 91989
rect 79619 91961 79647 91989
rect 79681 91961 79709 91989
rect 79743 91961 79771 91989
rect 79557 83147 79585 83175
rect 79619 83147 79647 83175
rect 79681 83147 79709 83175
rect 79743 83147 79771 83175
rect 79557 83085 79585 83113
rect 79619 83085 79647 83113
rect 79681 83085 79709 83113
rect 79743 83085 79771 83113
rect 79557 83023 79585 83051
rect 79619 83023 79647 83051
rect 79681 83023 79709 83051
rect 79743 83023 79771 83051
rect 79557 82961 79585 82989
rect 79619 82961 79647 82989
rect 79681 82961 79709 82989
rect 79743 82961 79771 82989
rect 79557 74147 79585 74175
rect 79619 74147 79647 74175
rect 79681 74147 79709 74175
rect 79743 74147 79771 74175
rect 79557 74085 79585 74113
rect 79619 74085 79647 74113
rect 79681 74085 79709 74113
rect 79743 74085 79771 74113
rect 79557 74023 79585 74051
rect 79619 74023 79647 74051
rect 79681 74023 79709 74051
rect 79743 74023 79771 74051
rect 79557 73961 79585 73989
rect 79619 73961 79647 73989
rect 79681 73961 79709 73989
rect 79743 73961 79771 73989
rect 79557 65147 79585 65175
rect 79619 65147 79647 65175
rect 79681 65147 79709 65175
rect 79743 65147 79771 65175
rect 79557 65085 79585 65113
rect 79619 65085 79647 65113
rect 79681 65085 79709 65113
rect 79743 65085 79771 65113
rect 79557 65023 79585 65051
rect 79619 65023 79647 65051
rect 79681 65023 79709 65051
rect 79743 65023 79771 65051
rect 79557 64961 79585 64989
rect 79619 64961 79647 64989
rect 79681 64961 79709 64989
rect 79743 64961 79771 64989
rect 79557 56147 79585 56175
rect 79619 56147 79647 56175
rect 79681 56147 79709 56175
rect 79743 56147 79771 56175
rect 79557 56085 79585 56113
rect 79619 56085 79647 56113
rect 79681 56085 79709 56113
rect 79743 56085 79771 56113
rect 79557 56023 79585 56051
rect 79619 56023 79647 56051
rect 79681 56023 79709 56051
rect 79743 56023 79771 56051
rect 79557 55961 79585 55989
rect 79619 55961 79647 55989
rect 79681 55961 79709 55989
rect 79743 55961 79771 55989
rect 79557 47147 79585 47175
rect 79619 47147 79647 47175
rect 79681 47147 79709 47175
rect 79743 47147 79771 47175
rect 79557 47085 79585 47113
rect 79619 47085 79647 47113
rect 79681 47085 79709 47113
rect 79743 47085 79771 47113
rect 79557 47023 79585 47051
rect 79619 47023 79647 47051
rect 79681 47023 79709 47051
rect 79743 47023 79771 47051
rect 79557 46961 79585 46989
rect 79619 46961 79647 46989
rect 79681 46961 79709 46989
rect 79743 46961 79771 46989
rect 79557 38147 79585 38175
rect 79619 38147 79647 38175
rect 79681 38147 79709 38175
rect 79743 38147 79771 38175
rect 79557 38085 79585 38113
rect 79619 38085 79647 38113
rect 79681 38085 79709 38113
rect 79743 38085 79771 38113
rect 79557 38023 79585 38051
rect 79619 38023 79647 38051
rect 79681 38023 79709 38051
rect 79743 38023 79771 38051
rect 79557 37961 79585 37989
rect 79619 37961 79647 37989
rect 79681 37961 79709 37989
rect 79743 37961 79771 37989
rect 79557 29147 79585 29175
rect 79619 29147 79647 29175
rect 79681 29147 79709 29175
rect 79743 29147 79771 29175
rect 79557 29085 79585 29113
rect 79619 29085 79647 29113
rect 79681 29085 79709 29113
rect 79743 29085 79771 29113
rect 79557 29023 79585 29051
rect 79619 29023 79647 29051
rect 79681 29023 79709 29051
rect 79743 29023 79771 29051
rect 79557 28961 79585 28989
rect 79619 28961 79647 28989
rect 79681 28961 79709 28989
rect 79743 28961 79771 28989
rect 79557 20147 79585 20175
rect 79619 20147 79647 20175
rect 79681 20147 79709 20175
rect 79743 20147 79771 20175
rect 79557 20085 79585 20113
rect 79619 20085 79647 20113
rect 79681 20085 79709 20113
rect 79743 20085 79771 20113
rect 79557 20023 79585 20051
rect 79619 20023 79647 20051
rect 79681 20023 79709 20051
rect 79743 20023 79771 20051
rect 79557 19961 79585 19989
rect 79619 19961 79647 19989
rect 79681 19961 79709 19989
rect 79743 19961 79771 19989
rect 79557 11147 79585 11175
rect 79619 11147 79647 11175
rect 79681 11147 79709 11175
rect 79743 11147 79771 11175
rect 79557 11085 79585 11113
rect 79619 11085 79647 11113
rect 79681 11085 79709 11113
rect 79743 11085 79771 11113
rect 79557 11023 79585 11051
rect 79619 11023 79647 11051
rect 79681 11023 79709 11051
rect 79743 11023 79771 11051
rect 79557 10961 79585 10989
rect 79619 10961 79647 10989
rect 79681 10961 79709 10989
rect 79743 10961 79771 10989
rect 79557 2147 79585 2175
rect 79619 2147 79647 2175
rect 79681 2147 79709 2175
rect 79743 2147 79771 2175
rect 79557 2085 79585 2113
rect 79619 2085 79647 2113
rect 79681 2085 79709 2113
rect 79743 2085 79771 2113
rect 79557 2023 79585 2051
rect 79619 2023 79647 2051
rect 79681 2023 79709 2051
rect 79743 2023 79771 2051
rect 79557 1961 79585 1989
rect 79619 1961 79647 1989
rect 79681 1961 79709 1989
rect 79743 1961 79771 1989
rect 79557 -108 79585 -80
rect 79619 -108 79647 -80
rect 79681 -108 79709 -80
rect 79743 -108 79771 -80
rect 79557 -170 79585 -142
rect 79619 -170 79647 -142
rect 79681 -170 79709 -142
rect 79743 -170 79771 -142
rect 79557 -232 79585 -204
rect 79619 -232 79647 -204
rect 79681 -232 79709 -204
rect 79743 -232 79771 -204
rect 79557 -294 79585 -266
rect 79619 -294 79647 -266
rect 79681 -294 79709 -266
rect 79743 -294 79771 -266
rect 81417 299058 81445 299086
rect 81479 299058 81507 299086
rect 81541 299058 81569 299086
rect 81603 299058 81631 299086
rect 81417 298996 81445 299024
rect 81479 298996 81507 299024
rect 81541 298996 81569 299024
rect 81603 298996 81631 299024
rect 81417 298934 81445 298962
rect 81479 298934 81507 298962
rect 81541 298934 81569 298962
rect 81603 298934 81631 298962
rect 81417 298872 81445 298900
rect 81479 298872 81507 298900
rect 81541 298872 81569 298900
rect 81603 298872 81631 298900
rect 81417 293147 81445 293175
rect 81479 293147 81507 293175
rect 81541 293147 81569 293175
rect 81603 293147 81631 293175
rect 81417 293085 81445 293113
rect 81479 293085 81507 293113
rect 81541 293085 81569 293113
rect 81603 293085 81631 293113
rect 81417 293023 81445 293051
rect 81479 293023 81507 293051
rect 81541 293023 81569 293051
rect 81603 293023 81631 293051
rect 81417 292961 81445 292989
rect 81479 292961 81507 292989
rect 81541 292961 81569 292989
rect 81603 292961 81631 292989
rect 81417 284147 81445 284175
rect 81479 284147 81507 284175
rect 81541 284147 81569 284175
rect 81603 284147 81631 284175
rect 81417 284085 81445 284113
rect 81479 284085 81507 284113
rect 81541 284085 81569 284113
rect 81603 284085 81631 284113
rect 81417 284023 81445 284051
rect 81479 284023 81507 284051
rect 81541 284023 81569 284051
rect 81603 284023 81631 284051
rect 81417 283961 81445 283989
rect 81479 283961 81507 283989
rect 81541 283961 81569 283989
rect 81603 283961 81631 283989
rect 81417 275147 81445 275175
rect 81479 275147 81507 275175
rect 81541 275147 81569 275175
rect 81603 275147 81631 275175
rect 81417 275085 81445 275113
rect 81479 275085 81507 275113
rect 81541 275085 81569 275113
rect 81603 275085 81631 275113
rect 81417 275023 81445 275051
rect 81479 275023 81507 275051
rect 81541 275023 81569 275051
rect 81603 275023 81631 275051
rect 81417 274961 81445 274989
rect 81479 274961 81507 274989
rect 81541 274961 81569 274989
rect 81603 274961 81631 274989
rect 81417 266147 81445 266175
rect 81479 266147 81507 266175
rect 81541 266147 81569 266175
rect 81603 266147 81631 266175
rect 81417 266085 81445 266113
rect 81479 266085 81507 266113
rect 81541 266085 81569 266113
rect 81603 266085 81631 266113
rect 81417 266023 81445 266051
rect 81479 266023 81507 266051
rect 81541 266023 81569 266051
rect 81603 266023 81631 266051
rect 81417 265961 81445 265989
rect 81479 265961 81507 265989
rect 81541 265961 81569 265989
rect 81603 265961 81631 265989
rect 81417 257147 81445 257175
rect 81479 257147 81507 257175
rect 81541 257147 81569 257175
rect 81603 257147 81631 257175
rect 81417 257085 81445 257113
rect 81479 257085 81507 257113
rect 81541 257085 81569 257113
rect 81603 257085 81631 257113
rect 81417 257023 81445 257051
rect 81479 257023 81507 257051
rect 81541 257023 81569 257051
rect 81603 257023 81631 257051
rect 81417 256961 81445 256989
rect 81479 256961 81507 256989
rect 81541 256961 81569 256989
rect 81603 256961 81631 256989
rect 81417 248147 81445 248175
rect 81479 248147 81507 248175
rect 81541 248147 81569 248175
rect 81603 248147 81631 248175
rect 81417 248085 81445 248113
rect 81479 248085 81507 248113
rect 81541 248085 81569 248113
rect 81603 248085 81631 248113
rect 81417 248023 81445 248051
rect 81479 248023 81507 248051
rect 81541 248023 81569 248051
rect 81603 248023 81631 248051
rect 81417 247961 81445 247989
rect 81479 247961 81507 247989
rect 81541 247961 81569 247989
rect 81603 247961 81631 247989
rect 81417 239147 81445 239175
rect 81479 239147 81507 239175
rect 81541 239147 81569 239175
rect 81603 239147 81631 239175
rect 81417 239085 81445 239113
rect 81479 239085 81507 239113
rect 81541 239085 81569 239113
rect 81603 239085 81631 239113
rect 81417 239023 81445 239051
rect 81479 239023 81507 239051
rect 81541 239023 81569 239051
rect 81603 239023 81631 239051
rect 81417 238961 81445 238989
rect 81479 238961 81507 238989
rect 81541 238961 81569 238989
rect 81603 238961 81631 238989
rect 81417 230147 81445 230175
rect 81479 230147 81507 230175
rect 81541 230147 81569 230175
rect 81603 230147 81631 230175
rect 81417 230085 81445 230113
rect 81479 230085 81507 230113
rect 81541 230085 81569 230113
rect 81603 230085 81631 230113
rect 81417 230023 81445 230051
rect 81479 230023 81507 230051
rect 81541 230023 81569 230051
rect 81603 230023 81631 230051
rect 81417 229961 81445 229989
rect 81479 229961 81507 229989
rect 81541 229961 81569 229989
rect 81603 229961 81631 229989
rect 81417 221147 81445 221175
rect 81479 221147 81507 221175
rect 81541 221147 81569 221175
rect 81603 221147 81631 221175
rect 81417 221085 81445 221113
rect 81479 221085 81507 221113
rect 81541 221085 81569 221113
rect 81603 221085 81631 221113
rect 81417 221023 81445 221051
rect 81479 221023 81507 221051
rect 81541 221023 81569 221051
rect 81603 221023 81631 221051
rect 81417 220961 81445 220989
rect 81479 220961 81507 220989
rect 81541 220961 81569 220989
rect 81603 220961 81631 220989
rect 81417 212147 81445 212175
rect 81479 212147 81507 212175
rect 81541 212147 81569 212175
rect 81603 212147 81631 212175
rect 81417 212085 81445 212113
rect 81479 212085 81507 212113
rect 81541 212085 81569 212113
rect 81603 212085 81631 212113
rect 81417 212023 81445 212051
rect 81479 212023 81507 212051
rect 81541 212023 81569 212051
rect 81603 212023 81631 212051
rect 81417 211961 81445 211989
rect 81479 211961 81507 211989
rect 81541 211961 81569 211989
rect 81603 211961 81631 211989
rect 81417 203147 81445 203175
rect 81479 203147 81507 203175
rect 81541 203147 81569 203175
rect 81603 203147 81631 203175
rect 81417 203085 81445 203113
rect 81479 203085 81507 203113
rect 81541 203085 81569 203113
rect 81603 203085 81631 203113
rect 81417 203023 81445 203051
rect 81479 203023 81507 203051
rect 81541 203023 81569 203051
rect 81603 203023 81631 203051
rect 81417 202961 81445 202989
rect 81479 202961 81507 202989
rect 81541 202961 81569 202989
rect 81603 202961 81631 202989
rect 81417 194147 81445 194175
rect 81479 194147 81507 194175
rect 81541 194147 81569 194175
rect 81603 194147 81631 194175
rect 81417 194085 81445 194113
rect 81479 194085 81507 194113
rect 81541 194085 81569 194113
rect 81603 194085 81631 194113
rect 81417 194023 81445 194051
rect 81479 194023 81507 194051
rect 81541 194023 81569 194051
rect 81603 194023 81631 194051
rect 81417 193961 81445 193989
rect 81479 193961 81507 193989
rect 81541 193961 81569 193989
rect 81603 193961 81631 193989
rect 81417 185147 81445 185175
rect 81479 185147 81507 185175
rect 81541 185147 81569 185175
rect 81603 185147 81631 185175
rect 81417 185085 81445 185113
rect 81479 185085 81507 185113
rect 81541 185085 81569 185113
rect 81603 185085 81631 185113
rect 81417 185023 81445 185051
rect 81479 185023 81507 185051
rect 81541 185023 81569 185051
rect 81603 185023 81631 185051
rect 81417 184961 81445 184989
rect 81479 184961 81507 184989
rect 81541 184961 81569 184989
rect 81603 184961 81631 184989
rect 81417 176147 81445 176175
rect 81479 176147 81507 176175
rect 81541 176147 81569 176175
rect 81603 176147 81631 176175
rect 81417 176085 81445 176113
rect 81479 176085 81507 176113
rect 81541 176085 81569 176113
rect 81603 176085 81631 176113
rect 81417 176023 81445 176051
rect 81479 176023 81507 176051
rect 81541 176023 81569 176051
rect 81603 176023 81631 176051
rect 81417 175961 81445 175989
rect 81479 175961 81507 175989
rect 81541 175961 81569 175989
rect 81603 175961 81631 175989
rect 81417 167147 81445 167175
rect 81479 167147 81507 167175
rect 81541 167147 81569 167175
rect 81603 167147 81631 167175
rect 81417 167085 81445 167113
rect 81479 167085 81507 167113
rect 81541 167085 81569 167113
rect 81603 167085 81631 167113
rect 81417 167023 81445 167051
rect 81479 167023 81507 167051
rect 81541 167023 81569 167051
rect 81603 167023 81631 167051
rect 81417 166961 81445 166989
rect 81479 166961 81507 166989
rect 81541 166961 81569 166989
rect 81603 166961 81631 166989
rect 81417 158147 81445 158175
rect 81479 158147 81507 158175
rect 81541 158147 81569 158175
rect 81603 158147 81631 158175
rect 81417 158085 81445 158113
rect 81479 158085 81507 158113
rect 81541 158085 81569 158113
rect 81603 158085 81631 158113
rect 81417 158023 81445 158051
rect 81479 158023 81507 158051
rect 81541 158023 81569 158051
rect 81603 158023 81631 158051
rect 81417 157961 81445 157989
rect 81479 157961 81507 157989
rect 81541 157961 81569 157989
rect 81603 157961 81631 157989
rect 81417 149147 81445 149175
rect 81479 149147 81507 149175
rect 81541 149147 81569 149175
rect 81603 149147 81631 149175
rect 81417 149085 81445 149113
rect 81479 149085 81507 149113
rect 81541 149085 81569 149113
rect 81603 149085 81631 149113
rect 81417 149023 81445 149051
rect 81479 149023 81507 149051
rect 81541 149023 81569 149051
rect 81603 149023 81631 149051
rect 81417 148961 81445 148989
rect 81479 148961 81507 148989
rect 81541 148961 81569 148989
rect 81603 148961 81631 148989
rect 81417 140147 81445 140175
rect 81479 140147 81507 140175
rect 81541 140147 81569 140175
rect 81603 140147 81631 140175
rect 81417 140085 81445 140113
rect 81479 140085 81507 140113
rect 81541 140085 81569 140113
rect 81603 140085 81631 140113
rect 81417 140023 81445 140051
rect 81479 140023 81507 140051
rect 81541 140023 81569 140051
rect 81603 140023 81631 140051
rect 81417 139961 81445 139989
rect 81479 139961 81507 139989
rect 81541 139961 81569 139989
rect 81603 139961 81631 139989
rect 81417 131147 81445 131175
rect 81479 131147 81507 131175
rect 81541 131147 81569 131175
rect 81603 131147 81631 131175
rect 81417 131085 81445 131113
rect 81479 131085 81507 131113
rect 81541 131085 81569 131113
rect 81603 131085 81631 131113
rect 81417 131023 81445 131051
rect 81479 131023 81507 131051
rect 81541 131023 81569 131051
rect 81603 131023 81631 131051
rect 81417 130961 81445 130989
rect 81479 130961 81507 130989
rect 81541 130961 81569 130989
rect 81603 130961 81631 130989
rect 81417 122147 81445 122175
rect 81479 122147 81507 122175
rect 81541 122147 81569 122175
rect 81603 122147 81631 122175
rect 81417 122085 81445 122113
rect 81479 122085 81507 122113
rect 81541 122085 81569 122113
rect 81603 122085 81631 122113
rect 81417 122023 81445 122051
rect 81479 122023 81507 122051
rect 81541 122023 81569 122051
rect 81603 122023 81631 122051
rect 81417 121961 81445 121989
rect 81479 121961 81507 121989
rect 81541 121961 81569 121989
rect 81603 121961 81631 121989
rect 81417 113147 81445 113175
rect 81479 113147 81507 113175
rect 81541 113147 81569 113175
rect 81603 113147 81631 113175
rect 81417 113085 81445 113113
rect 81479 113085 81507 113113
rect 81541 113085 81569 113113
rect 81603 113085 81631 113113
rect 81417 113023 81445 113051
rect 81479 113023 81507 113051
rect 81541 113023 81569 113051
rect 81603 113023 81631 113051
rect 81417 112961 81445 112989
rect 81479 112961 81507 112989
rect 81541 112961 81569 112989
rect 81603 112961 81631 112989
rect 81417 104147 81445 104175
rect 81479 104147 81507 104175
rect 81541 104147 81569 104175
rect 81603 104147 81631 104175
rect 81417 104085 81445 104113
rect 81479 104085 81507 104113
rect 81541 104085 81569 104113
rect 81603 104085 81631 104113
rect 81417 104023 81445 104051
rect 81479 104023 81507 104051
rect 81541 104023 81569 104051
rect 81603 104023 81631 104051
rect 81417 103961 81445 103989
rect 81479 103961 81507 103989
rect 81541 103961 81569 103989
rect 81603 103961 81631 103989
rect 81417 95147 81445 95175
rect 81479 95147 81507 95175
rect 81541 95147 81569 95175
rect 81603 95147 81631 95175
rect 81417 95085 81445 95113
rect 81479 95085 81507 95113
rect 81541 95085 81569 95113
rect 81603 95085 81631 95113
rect 81417 95023 81445 95051
rect 81479 95023 81507 95051
rect 81541 95023 81569 95051
rect 81603 95023 81631 95051
rect 81417 94961 81445 94989
rect 81479 94961 81507 94989
rect 81541 94961 81569 94989
rect 81603 94961 81631 94989
rect 81417 86147 81445 86175
rect 81479 86147 81507 86175
rect 81541 86147 81569 86175
rect 81603 86147 81631 86175
rect 81417 86085 81445 86113
rect 81479 86085 81507 86113
rect 81541 86085 81569 86113
rect 81603 86085 81631 86113
rect 81417 86023 81445 86051
rect 81479 86023 81507 86051
rect 81541 86023 81569 86051
rect 81603 86023 81631 86051
rect 81417 85961 81445 85989
rect 81479 85961 81507 85989
rect 81541 85961 81569 85989
rect 81603 85961 81631 85989
rect 81417 77147 81445 77175
rect 81479 77147 81507 77175
rect 81541 77147 81569 77175
rect 81603 77147 81631 77175
rect 81417 77085 81445 77113
rect 81479 77085 81507 77113
rect 81541 77085 81569 77113
rect 81603 77085 81631 77113
rect 81417 77023 81445 77051
rect 81479 77023 81507 77051
rect 81541 77023 81569 77051
rect 81603 77023 81631 77051
rect 81417 76961 81445 76989
rect 81479 76961 81507 76989
rect 81541 76961 81569 76989
rect 81603 76961 81631 76989
rect 81417 68147 81445 68175
rect 81479 68147 81507 68175
rect 81541 68147 81569 68175
rect 81603 68147 81631 68175
rect 81417 68085 81445 68113
rect 81479 68085 81507 68113
rect 81541 68085 81569 68113
rect 81603 68085 81631 68113
rect 81417 68023 81445 68051
rect 81479 68023 81507 68051
rect 81541 68023 81569 68051
rect 81603 68023 81631 68051
rect 81417 67961 81445 67989
rect 81479 67961 81507 67989
rect 81541 67961 81569 67989
rect 81603 67961 81631 67989
rect 81417 59147 81445 59175
rect 81479 59147 81507 59175
rect 81541 59147 81569 59175
rect 81603 59147 81631 59175
rect 81417 59085 81445 59113
rect 81479 59085 81507 59113
rect 81541 59085 81569 59113
rect 81603 59085 81631 59113
rect 81417 59023 81445 59051
rect 81479 59023 81507 59051
rect 81541 59023 81569 59051
rect 81603 59023 81631 59051
rect 81417 58961 81445 58989
rect 81479 58961 81507 58989
rect 81541 58961 81569 58989
rect 81603 58961 81631 58989
rect 81417 50147 81445 50175
rect 81479 50147 81507 50175
rect 81541 50147 81569 50175
rect 81603 50147 81631 50175
rect 81417 50085 81445 50113
rect 81479 50085 81507 50113
rect 81541 50085 81569 50113
rect 81603 50085 81631 50113
rect 81417 50023 81445 50051
rect 81479 50023 81507 50051
rect 81541 50023 81569 50051
rect 81603 50023 81631 50051
rect 81417 49961 81445 49989
rect 81479 49961 81507 49989
rect 81541 49961 81569 49989
rect 81603 49961 81631 49989
rect 81417 41147 81445 41175
rect 81479 41147 81507 41175
rect 81541 41147 81569 41175
rect 81603 41147 81631 41175
rect 81417 41085 81445 41113
rect 81479 41085 81507 41113
rect 81541 41085 81569 41113
rect 81603 41085 81631 41113
rect 81417 41023 81445 41051
rect 81479 41023 81507 41051
rect 81541 41023 81569 41051
rect 81603 41023 81631 41051
rect 81417 40961 81445 40989
rect 81479 40961 81507 40989
rect 81541 40961 81569 40989
rect 81603 40961 81631 40989
rect 81417 32147 81445 32175
rect 81479 32147 81507 32175
rect 81541 32147 81569 32175
rect 81603 32147 81631 32175
rect 81417 32085 81445 32113
rect 81479 32085 81507 32113
rect 81541 32085 81569 32113
rect 81603 32085 81631 32113
rect 81417 32023 81445 32051
rect 81479 32023 81507 32051
rect 81541 32023 81569 32051
rect 81603 32023 81631 32051
rect 81417 31961 81445 31989
rect 81479 31961 81507 31989
rect 81541 31961 81569 31989
rect 81603 31961 81631 31989
rect 81417 23147 81445 23175
rect 81479 23147 81507 23175
rect 81541 23147 81569 23175
rect 81603 23147 81631 23175
rect 81417 23085 81445 23113
rect 81479 23085 81507 23113
rect 81541 23085 81569 23113
rect 81603 23085 81631 23113
rect 81417 23023 81445 23051
rect 81479 23023 81507 23051
rect 81541 23023 81569 23051
rect 81603 23023 81631 23051
rect 81417 22961 81445 22989
rect 81479 22961 81507 22989
rect 81541 22961 81569 22989
rect 81603 22961 81631 22989
rect 81417 14147 81445 14175
rect 81479 14147 81507 14175
rect 81541 14147 81569 14175
rect 81603 14147 81631 14175
rect 81417 14085 81445 14113
rect 81479 14085 81507 14113
rect 81541 14085 81569 14113
rect 81603 14085 81631 14113
rect 81417 14023 81445 14051
rect 81479 14023 81507 14051
rect 81541 14023 81569 14051
rect 81603 14023 81631 14051
rect 81417 13961 81445 13989
rect 81479 13961 81507 13989
rect 81541 13961 81569 13989
rect 81603 13961 81631 13989
rect 81417 5147 81445 5175
rect 81479 5147 81507 5175
rect 81541 5147 81569 5175
rect 81603 5147 81631 5175
rect 81417 5085 81445 5113
rect 81479 5085 81507 5113
rect 81541 5085 81569 5113
rect 81603 5085 81631 5113
rect 81417 5023 81445 5051
rect 81479 5023 81507 5051
rect 81541 5023 81569 5051
rect 81603 5023 81631 5051
rect 81417 4961 81445 4989
rect 81479 4961 81507 4989
rect 81541 4961 81569 4989
rect 81603 4961 81631 4989
rect 81417 -588 81445 -560
rect 81479 -588 81507 -560
rect 81541 -588 81569 -560
rect 81603 -588 81631 -560
rect 81417 -650 81445 -622
rect 81479 -650 81507 -622
rect 81541 -650 81569 -622
rect 81603 -650 81631 -622
rect 81417 -712 81445 -684
rect 81479 -712 81507 -684
rect 81541 -712 81569 -684
rect 81603 -712 81631 -684
rect 81417 -774 81445 -746
rect 81479 -774 81507 -746
rect 81541 -774 81569 -746
rect 81603 -774 81631 -746
rect 94917 298578 94945 298606
rect 94979 298578 95007 298606
rect 95041 298578 95069 298606
rect 95103 298578 95131 298606
rect 94917 298516 94945 298544
rect 94979 298516 95007 298544
rect 95041 298516 95069 298544
rect 95103 298516 95131 298544
rect 94917 298454 94945 298482
rect 94979 298454 95007 298482
rect 95041 298454 95069 298482
rect 95103 298454 95131 298482
rect 94917 298392 94945 298420
rect 94979 298392 95007 298420
rect 95041 298392 95069 298420
rect 95103 298392 95131 298420
rect 94917 290147 94945 290175
rect 94979 290147 95007 290175
rect 95041 290147 95069 290175
rect 95103 290147 95131 290175
rect 94917 290085 94945 290113
rect 94979 290085 95007 290113
rect 95041 290085 95069 290113
rect 95103 290085 95131 290113
rect 94917 290023 94945 290051
rect 94979 290023 95007 290051
rect 95041 290023 95069 290051
rect 95103 290023 95131 290051
rect 94917 289961 94945 289989
rect 94979 289961 95007 289989
rect 95041 289961 95069 289989
rect 95103 289961 95131 289989
rect 94917 281147 94945 281175
rect 94979 281147 95007 281175
rect 95041 281147 95069 281175
rect 95103 281147 95131 281175
rect 94917 281085 94945 281113
rect 94979 281085 95007 281113
rect 95041 281085 95069 281113
rect 95103 281085 95131 281113
rect 94917 281023 94945 281051
rect 94979 281023 95007 281051
rect 95041 281023 95069 281051
rect 95103 281023 95131 281051
rect 94917 280961 94945 280989
rect 94979 280961 95007 280989
rect 95041 280961 95069 280989
rect 95103 280961 95131 280989
rect 94917 272147 94945 272175
rect 94979 272147 95007 272175
rect 95041 272147 95069 272175
rect 95103 272147 95131 272175
rect 94917 272085 94945 272113
rect 94979 272085 95007 272113
rect 95041 272085 95069 272113
rect 95103 272085 95131 272113
rect 94917 272023 94945 272051
rect 94979 272023 95007 272051
rect 95041 272023 95069 272051
rect 95103 272023 95131 272051
rect 94917 271961 94945 271989
rect 94979 271961 95007 271989
rect 95041 271961 95069 271989
rect 95103 271961 95131 271989
rect 94917 263147 94945 263175
rect 94979 263147 95007 263175
rect 95041 263147 95069 263175
rect 95103 263147 95131 263175
rect 94917 263085 94945 263113
rect 94979 263085 95007 263113
rect 95041 263085 95069 263113
rect 95103 263085 95131 263113
rect 94917 263023 94945 263051
rect 94979 263023 95007 263051
rect 95041 263023 95069 263051
rect 95103 263023 95131 263051
rect 94917 262961 94945 262989
rect 94979 262961 95007 262989
rect 95041 262961 95069 262989
rect 95103 262961 95131 262989
rect 94917 254147 94945 254175
rect 94979 254147 95007 254175
rect 95041 254147 95069 254175
rect 95103 254147 95131 254175
rect 94917 254085 94945 254113
rect 94979 254085 95007 254113
rect 95041 254085 95069 254113
rect 95103 254085 95131 254113
rect 94917 254023 94945 254051
rect 94979 254023 95007 254051
rect 95041 254023 95069 254051
rect 95103 254023 95131 254051
rect 94917 253961 94945 253989
rect 94979 253961 95007 253989
rect 95041 253961 95069 253989
rect 95103 253961 95131 253989
rect 94917 245147 94945 245175
rect 94979 245147 95007 245175
rect 95041 245147 95069 245175
rect 95103 245147 95131 245175
rect 94917 245085 94945 245113
rect 94979 245085 95007 245113
rect 95041 245085 95069 245113
rect 95103 245085 95131 245113
rect 94917 245023 94945 245051
rect 94979 245023 95007 245051
rect 95041 245023 95069 245051
rect 95103 245023 95131 245051
rect 94917 244961 94945 244989
rect 94979 244961 95007 244989
rect 95041 244961 95069 244989
rect 95103 244961 95131 244989
rect 94917 236147 94945 236175
rect 94979 236147 95007 236175
rect 95041 236147 95069 236175
rect 95103 236147 95131 236175
rect 94917 236085 94945 236113
rect 94979 236085 95007 236113
rect 95041 236085 95069 236113
rect 95103 236085 95131 236113
rect 94917 236023 94945 236051
rect 94979 236023 95007 236051
rect 95041 236023 95069 236051
rect 95103 236023 95131 236051
rect 94917 235961 94945 235989
rect 94979 235961 95007 235989
rect 95041 235961 95069 235989
rect 95103 235961 95131 235989
rect 94917 227147 94945 227175
rect 94979 227147 95007 227175
rect 95041 227147 95069 227175
rect 95103 227147 95131 227175
rect 94917 227085 94945 227113
rect 94979 227085 95007 227113
rect 95041 227085 95069 227113
rect 95103 227085 95131 227113
rect 94917 227023 94945 227051
rect 94979 227023 95007 227051
rect 95041 227023 95069 227051
rect 95103 227023 95131 227051
rect 94917 226961 94945 226989
rect 94979 226961 95007 226989
rect 95041 226961 95069 226989
rect 95103 226961 95131 226989
rect 94917 218147 94945 218175
rect 94979 218147 95007 218175
rect 95041 218147 95069 218175
rect 95103 218147 95131 218175
rect 94917 218085 94945 218113
rect 94979 218085 95007 218113
rect 95041 218085 95069 218113
rect 95103 218085 95131 218113
rect 94917 218023 94945 218051
rect 94979 218023 95007 218051
rect 95041 218023 95069 218051
rect 95103 218023 95131 218051
rect 94917 217961 94945 217989
rect 94979 217961 95007 217989
rect 95041 217961 95069 217989
rect 95103 217961 95131 217989
rect 94917 209147 94945 209175
rect 94979 209147 95007 209175
rect 95041 209147 95069 209175
rect 95103 209147 95131 209175
rect 94917 209085 94945 209113
rect 94979 209085 95007 209113
rect 95041 209085 95069 209113
rect 95103 209085 95131 209113
rect 94917 209023 94945 209051
rect 94979 209023 95007 209051
rect 95041 209023 95069 209051
rect 95103 209023 95131 209051
rect 94917 208961 94945 208989
rect 94979 208961 95007 208989
rect 95041 208961 95069 208989
rect 95103 208961 95131 208989
rect 94917 200147 94945 200175
rect 94979 200147 95007 200175
rect 95041 200147 95069 200175
rect 95103 200147 95131 200175
rect 94917 200085 94945 200113
rect 94979 200085 95007 200113
rect 95041 200085 95069 200113
rect 95103 200085 95131 200113
rect 94917 200023 94945 200051
rect 94979 200023 95007 200051
rect 95041 200023 95069 200051
rect 95103 200023 95131 200051
rect 94917 199961 94945 199989
rect 94979 199961 95007 199989
rect 95041 199961 95069 199989
rect 95103 199961 95131 199989
rect 94917 191147 94945 191175
rect 94979 191147 95007 191175
rect 95041 191147 95069 191175
rect 95103 191147 95131 191175
rect 94917 191085 94945 191113
rect 94979 191085 95007 191113
rect 95041 191085 95069 191113
rect 95103 191085 95131 191113
rect 94917 191023 94945 191051
rect 94979 191023 95007 191051
rect 95041 191023 95069 191051
rect 95103 191023 95131 191051
rect 94917 190961 94945 190989
rect 94979 190961 95007 190989
rect 95041 190961 95069 190989
rect 95103 190961 95131 190989
rect 94917 182147 94945 182175
rect 94979 182147 95007 182175
rect 95041 182147 95069 182175
rect 95103 182147 95131 182175
rect 94917 182085 94945 182113
rect 94979 182085 95007 182113
rect 95041 182085 95069 182113
rect 95103 182085 95131 182113
rect 94917 182023 94945 182051
rect 94979 182023 95007 182051
rect 95041 182023 95069 182051
rect 95103 182023 95131 182051
rect 94917 181961 94945 181989
rect 94979 181961 95007 181989
rect 95041 181961 95069 181989
rect 95103 181961 95131 181989
rect 94917 173147 94945 173175
rect 94979 173147 95007 173175
rect 95041 173147 95069 173175
rect 95103 173147 95131 173175
rect 94917 173085 94945 173113
rect 94979 173085 95007 173113
rect 95041 173085 95069 173113
rect 95103 173085 95131 173113
rect 94917 173023 94945 173051
rect 94979 173023 95007 173051
rect 95041 173023 95069 173051
rect 95103 173023 95131 173051
rect 94917 172961 94945 172989
rect 94979 172961 95007 172989
rect 95041 172961 95069 172989
rect 95103 172961 95131 172989
rect 94917 164147 94945 164175
rect 94979 164147 95007 164175
rect 95041 164147 95069 164175
rect 95103 164147 95131 164175
rect 94917 164085 94945 164113
rect 94979 164085 95007 164113
rect 95041 164085 95069 164113
rect 95103 164085 95131 164113
rect 94917 164023 94945 164051
rect 94979 164023 95007 164051
rect 95041 164023 95069 164051
rect 95103 164023 95131 164051
rect 94917 163961 94945 163989
rect 94979 163961 95007 163989
rect 95041 163961 95069 163989
rect 95103 163961 95131 163989
rect 94917 155147 94945 155175
rect 94979 155147 95007 155175
rect 95041 155147 95069 155175
rect 95103 155147 95131 155175
rect 94917 155085 94945 155113
rect 94979 155085 95007 155113
rect 95041 155085 95069 155113
rect 95103 155085 95131 155113
rect 94917 155023 94945 155051
rect 94979 155023 95007 155051
rect 95041 155023 95069 155051
rect 95103 155023 95131 155051
rect 94917 154961 94945 154989
rect 94979 154961 95007 154989
rect 95041 154961 95069 154989
rect 95103 154961 95131 154989
rect 94917 146147 94945 146175
rect 94979 146147 95007 146175
rect 95041 146147 95069 146175
rect 95103 146147 95131 146175
rect 94917 146085 94945 146113
rect 94979 146085 95007 146113
rect 95041 146085 95069 146113
rect 95103 146085 95131 146113
rect 94917 146023 94945 146051
rect 94979 146023 95007 146051
rect 95041 146023 95069 146051
rect 95103 146023 95131 146051
rect 94917 145961 94945 145989
rect 94979 145961 95007 145989
rect 95041 145961 95069 145989
rect 95103 145961 95131 145989
rect 94917 137147 94945 137175
rect 94979 137147 95007 137175
rect 95041 137147 95069 137175
rect 95103 137147 95131 137175
rect 94917 137085 94945 137113
rect 94979 137085 95007 137113
rect 95041 137085 95069 137113
rect 95103 137085 95131 137113
rect 94917 137023 94945 137051
rect 94979 137023 95007 137051
rect 95041 137023 95069 137051
rect 95103 137023 95131 137051
rect 94917 136961 94945 136989
rect 94979 136961 95007 136989
rect 95041 136961 95069 136989
rect 95103 136961 95131 136989
rect 94917 128147 94945 128175
rect 94979 128147 95007 128175
rect 95041 128147 95069 128175
rect 95103 128147 95131 128175
rect 94917 128085 94945 128113
rect 94979 128085 95007 128113
rect 95041 128085 95069 128113
rect 95103 128085 95131 128113
rect 94917 128023 94945 128051
rect 94979 128023 95007 128051
rect 95041 128023 95069 128051
rect 95103 128023 95131 128051
rect 94917 127961 94945 127989
rect 94979 127961 95007 127989
rect 95041 127961 95069 127989
rect 95103 127961 95131 127989
rect 94917 119147 94945 119175
rect 94979 119147 95007 119175
rect 95041 119147 95069 119175
rect 95103 119147 95131 119175
rect 94917 119085 94945 119113
rect 94979 119085 95007 119113
rect 95041 119085 95069 119113
rect 95103 119085 95131 119113
rect 94917 119023 94945 119051
rect 94979 119023 95007 119051
rect 95041 119023 95069 119051
rect 95103 119023 95131 119051
rect 94917 118961 94945 118989
rect 94979 118961 95007 118989
rect 95041 118961 95069 118989
rect 95103 118961 95131 118989
rect 94917 110147 94945 110175
rect 94979 110147 95007 110175
rect 95041 110147 95069 110175
rect 95103 110147 95131 110175
rect 94917 110085 94945 110113
rect 94979 110085 95007 110113
rect 95041 110085 95069 110113
rect 95103 110085 95131 110113
rect 94917 110023 94945 110051
rect 94979 110023 95007 110051
rect 95041 110023 95069 110051
rect 95103 110023 95131 110051
rect 94917 109961 94945 109989
rect 94979 109961 95007 109989
rect 95041 109961 95069 109989
rect 95103 109961 95131 109989
rect 94917 101147 94945 101175
rect 94979 101147 95007 101175
rect 95041 101147 95069 101175
rect 95103 101147 95131 101175
rect 94917 101085 94945 101113
rect 94979 101085 95007 101113
rect 95041 101085 95069 101113
rect 95103 101085 95131 101113
rect 94917 101023 94945 101051
rect 94979 101023 95007 101051
rect 95041 101023 95069 101051
rect 95103 101023 95131 101051
rect 94917 100961 94945 100989
rect 94979 100961 95007 100989
rect 95041 100961 95069 100989
rect 95103 100961 95131 100989
rect 94917 92147 94945 92175
rect 94979 92147 95007 92175
rect 95041 92147 95069 92175
rect 95103 92147 95131 92175
rect 94917 92085 94945 92113
rect 94979 92085 95007 92113
rect 95041 92085 95069 92113
rect 95103 92085 95131 92113
rect 94917 92023 94945 92051
rect 94979 92023 95007 92051
rect 95041 92023 95069 92051
rect 95103 92023 95131 92051
rect 94917 91961 94945 91989
rect 94979 91961 95007 91989
rect 95041 91961 95069 91989
rect 95103 91961 95131 91989
rect 94917 83147 94945 83175
rect 94979 83147 95007 83175
rect 95041 83147 95069 83175
rect 95103 83147 95131 83175
rect 94917 83085 94945 83113
rect 94979 83085 95007 83113
rect 95041 83085 95069 83113
rect 95103 83085 95131 83113
rect 94917 83023 94945 83051
rect 94979 83023 95007 83051
rect 95041 83023 95069 83051
rect 95103 83023 95131 83051
rect 94917 82961 94945 82989
rect 94979 82961 95007 82989
rect 95041 82961 95069 82989
rect 95103 82961 95131 82989
rect 94917 74147 94945 74175
rect 94979 74147 95007 74175
rect 95041 74147 95069 74175
rect 95103 74147 95131 74175
rect 94917 74085 94945 74113
rect 94979 74085 95007 74113
rect 95041 74085 95069 74113
rect 95103 74085 95131 74113
rect 94917 74023 94945 74051
rect 94979 74023 95007 74051
rect 95041 74023 95069 74051
rect 95103 74023 95131 74051
rect 94917 73961 94945 73989
rect 94979 73961 95007 73989
rect 95041 73961 95069 73989
rect 95103 73961 95131 73989
rect 94917 65147 94945 65175
rect 94979 65147 95007 65175
rect 95041 65147 95069 65175
rect 95103 65147 95131 65175
rect 94917 65085 94945 65113
rect 94979 65085 95007 65113
rect 95041 65085 95069 65113
rect 95103 65085 95131 65113
rect 94917 65023 94945 65051
rect 94979 65023 95007 65051
rect 95041 65023 95069 65051
rect 95103 65023 95131 65051
rect 94917 64961 94945 64989
rect 94979 64961 95007 64989
rect 95041 64961 95069 64989
rect 95103 64961 95131 64989
rect 94917 56147 94945 56175
rect 94979 56147 95007 56175
rect 95041 56147 95069 56175
rect 95103 56147 95131 56175
rect 94917 56085 94945 56113
rect 94979 56085 95007 56113
rect 95041 56085 95069 56113
rect 95103 56085 95131 56113
rect 94917 56023 94945 56051
rect 94979 56023 95007 56051
rect 95041 56023 95069 56051
rect 95103 56023 95131 56051
rect 94917 55961 94945 55989
rect 94979 55961 95007 55989
rect 95041 55961 95069 55989
rect 95103 55961 95131 55989
rect 94917 47147 94945 47175
rect 94979 47147 95007 47175
rect 95041 47147 95069 47175
rect 95103 47147 95131 47175
rect 94917 47085 94945 47113
rect 94979 47085 95007 47113
rect 95041 47085 95069 47113
rect 95103 47085 95131 47113
rect 94917 47023 94945 47051
rect 94979 47023 95007 47051
rect 95041 47023 95069 47051
rect 95103 47023 95131 47051
rect 94917 46961 94945 46989
rect 94979 46961 95007 46989
rect 95041 46961 95069 46989
rect 95103 46961 95131 46989
rect 94917 38147 94945 38175
rect 94979 38147 95007 38175
rect 95041 38147 95069 38175
rect 95103 38147 95131 38175
rect 94917 38085 94945 38113
rect 94979 38085 95007 38113
rect 95041 38085 95069 38113
rect 95103 38085 95131 38113
rect 94917 38023 94945 38051
rect 94979 38023 95007 38051
rect 95041 38023 95069 38051
rect 95103 38023 95131 38051
rect 94917 37961 94945 37989
rect 94979 37961 95007 37989
rect 95041 37961 95069 37989
rect 95103 37961 95131 37989
rect 94917 29147 94945 29175
rect 94979 29147 95007 29175
rect 95041 29147 95069 29175
rect 95103 29147 95131 29175
rect 94917 29085 94945 29113
rect 94979 29085 95007 29113
rect 95041 29085 95069 29113
rect 95103 29085 95131 29113
rect 94917 29023 94945 29051
rect 94979 29023 95007 29051
rect 95041 29023 95069 29051
rect 95103 29023 95131 29051
rect 94917 28961 94945 28989
rect 94979 28961 95007 28989
rect 95041 28961 95069 28989
rect 95103 28961 95131 28989
rect 94917 20147 94945 20175
rect 94979 20147 95007 20175
rect 95041 20147 95069 20175
rect 95103 20147 95131 20175
rect 94917 20085 94945 20113
rect 94979 20085 95007 20113
rect 95041 20085 95069 20113
rect 95103 20085 95131 20113
rect 94917 20023 94945 20051
rect 94979 20023 95007 20051
rect 95041 20023 95069 20051
rect 95103 20023 95131 20051
rect 94917 19961 94945 19989
rect 94979 19961 95007 19989
rect 95041 19961 95069 19989
rect 95103 19961 95131 19989
rect 94917 11147 94945 11175
rect 94979 11147 95007 11175
rect 95041 11147 95069 11175
rect 95103 11147 95131 11175
rect 94917 11085 94945 11113
rect 94979 11085 95007 11113
rect 95041 11085 95069 11113
rect 95103 11085 95131 11113
rect 94917 11023 94945 11051
rect 94979 11023 95007 11051
rect 95041 11023 95069 11051
rect 95103 11023 95131 11051
rect 94917 10961 94945 10989
rect 94979 10961 95007 10989
rect 95041 10961 95069 10989
rect 95103 10961 95131 10989
rect 94917 2147 94945 2175
rect 94979 2147 95007 2175
rect 95041 2147 95069 2175
rect 95103 2147 95131 2175
rect 94917 2085 94945 2113
rect 94979 2085 95007 2113
rect 95041 2085 95069 2113
rect 95103 2085 95131 2113
rect 94917 2023 94945 2051
rect 94979 2023 95007 2051
rect 95041 2023 95069 2051
rect 95103 2023 95131 2051
rect 94917 1961 94945 1989
rect 94979 1961 95007 1989
rect 95041 1961 95069 1989
rect 95103 1961 95131 1989
rect 94917 -108 94945 -80
rect 94979 -108 95007 -80
rect 95041 -108 95069 -80
rect 95103 -108 95131 -80
rect 94917 -170 94945 -142
rect 94979 -170 95007 -142
rect 95041 -170 95069 -142
rect 95103 -170 95131 -142
rect 94917 -232 94945 -204
rect 94979 -232 95007 -204
rect 95041 -232 95069 -204
rect 95103 -232 95131 -204
rect 94917 -294 94945 -266
rect 94979 -294 95007 -266
rect 95041 -294 95069 -266
rect 95103 -294 95131 -266
rect 96777 299058 96805 299086
rect 96839 299058 96867 299086
rect 96901 299058 96929 299086
rect 96963 299058 96991 299086
rect 96777 298996 96805 299024
rect 96839 298996 96867 299024
rect 96901 298996 96929 299024
rect 96963 298996 96991 299024
rect 96777 298934 96805 298962
rect 96839 298934 96867 298962
rect 96901 298934 96929 298962
rect 96963 298934 96991 298962
rect 96777 298872 96805 298900
rect 96839 298872 96867 298900
rect 96901 298872 96929 298900
rect 96963 298872 96991 298900
rect 96777 293147 96805 293175
rect 96839 293147 96867 293175
rect 96901 293147 96929 293175
rect 96963 293147 96991 293175
rect 96777 293085 96805 293113
rect 96839 293085 96867 293113
rect 96901 293085 96929 293113
rect 96963 293085 96991 293113
rect 96777 293023 96805 293051
rect 96839 293023 96867 293051
rect 96901 293023 96929 293051
rect 96963 293023 96991 293051
rect 96777 292961 96805 292989
rect 96839 292961 96867 292989
rect 96901 292961 96929 292989
rect 96963 292961 96991 292989
rect 96777 284147 96805 284175
rect 96839 284147 96867 284175
rect 96901 284147 96929 284175
rect 96963 284147 96991 284175
rect 96777 284085 96805 284113
rect 96839 284085 96867 284113
rect 96901 284085 96929 284113
rect 96963 284085 96991 284113
rect 96777 284023 96805 284051
rect 96839 284023 96867 284051
rect 96901 284023 96929 284051
rect 96963 284023 96991 284051
rect 96777 283961 96805 283989
rect 96839 283961 96867 283989
rect 96901 283961 96929 283989
rect 96963 283961 96991 283989
rect 110277 298578 110305 298606
rect 110339 298578 110367 298606
rect 110401 298578 110429 298606
rect 110463 298578 110491 298606
rect 110277 298516 110305 298544
rect 110339 298516 110367 298544
rect 110401 298516 110429 298544
rect 110463 298516 110491 298544
rect 110277 298454 110305 298482
rect 110339 298454 110367 298482
rect 110401 298454 110429 298482
rect 110463 298454 110491 298482
rect 110277 298392 110305 298420
rect 110339 298392 110367 298420
rect 110401 298392 110429 298420
rect 110463 298392 110491 298420
rect 110277 290147 110305 290175
rect 110339 290147 110367 290175
rect 110401 290147 110429 290175
rect 110463 290147 110491 290175
rect 110277 290085 110305 290113
rect 110339 290085 110367 290113
rect 110401 290085 110429 290113
rect 110463 290085 110491 290113
rect 110277 290023 110305 290051
rect 110339 290023 110367 290051
rect 110401 290023 110429 290051
rect 110463 290023 110491 290051
rect 110277 289961 110305 289989
rect 110339 289961 110367 289989
rect 110401 289961 110429 289989
rect 110463 289961 110491 289989
rect 110277 281147 110305 281175
rect 110339 281147 110367 281175
rect 110401 281147 110429 281175
rect 110463 281147 110491 281175
rect 110277 281085 110305 281113
rect 110339 281085 110367 281113
rect 110401 281085 110429 281113
rect 110463 281085 110491 281113
rect 110277 281023 110305 281051
rect 110339 281023 110367 281051
rect 110401 281023 110429 281051
rect 110463 281023 110491 281051
rect 110277 280961 110305 280989
rect 110339 280961 110367 280989
rect 110401 280961 110429 280989
rect 110463 280961 110491 280989
rect 112137 299058 112165 299086
rect 112199 299058 112227 299086
rect 112261 299058 112289 299086
rect 112323 299058 112351 299086
rect 112137 298996 112165 299024
rect 112199 298996 112227 299024
rect 112261 298996 112289 299024
rect 112323 298996 112351 299024
rect 112137 298934 112165 298962
rect 112199 298934 112227 298962
rect 112261 298934 112289 298962
rect 112323 298934 112351 298962
rect 112137 298872 112165 298900
rect 112199 298872 112227 298900
rect 112261 298872 112289 298900
rect 112323 298872 112351 298900
rect 112137 293147 112165 293175
rect 112199 293147 112227 293175
rect 112261 293147 112289 293175
rect 112323 293147 112351 293175
rect 112137 293085 112165 293113
rect 112199 293085 112227 293113
rect 112261 293085 112289 293113
rect 112323 293085 112351 293113
rect 112137 293023 112165 293051
rect 112199 293023 112227 293051
rect 112261 293023 112289 293051
rect 112323 293023 112351 293051
rect 112137 292961 112165 292989
rect 112199 292961 112227 292989
rect 112261 292961 112289 292989
rect 112323 292961 112351 292989
rect 112137 284147 112165 284175
rect 112199 284147 112227 284175
rect 112261 284147 112289 284175
rect 112323 284147 112351 284175
rect 112137 284085 112165 284113
rect 112199 284085 112227 284113
rect 112261 284085 112289 284113
rect 112323 284085 112351 284113
rect 112137 284023 112165 284051
rect 112199 284023 112227 284051
rect 112261 284023 112289 284051
rect 112323 284023 112351 284051
rect 112137 283961 112165 283989
rect 112199 283961 112227 283989
rect 112261 283961 112289 283989
rect 112323 283961 112351 283989
rect 125637 298578 125665 298606
rect 125699 298578 125727 298606
rect 125761 298578 125789 298606
rect 125823 298578 125851 298606
rect 125637 298516 125665 298544
rect 125699 298516 125727 298544
rect 125761 298516 125789 298544
rect 125823 298516 125851 298544
rect 125637 298454 125665 298482
rect 125699 298454 125727 298482
rect 125761 298454 125789 298482
rect 125823 298454 125851 298482
rect 125637 298392 125665 298420
rect 125699 298392 125727 298420
rect 125761 298392 125789 298420
rect 125823 298392 125851 298420
rect 125637 290147 125665 290175
rect 125699 290147 125727 290175
rect 125761 290147 125789 290175
rect 125823 290147 125851 290175
rect 125637 290085 125665 290113
rect 125699 290085 125727 290113
rect 125761 290085 125789 290113
rect 125823 290085 125851 290113
rect 125637 290023 125665 290051
rect 125699 290023 125727 290051
rect 125761 290023 125789 290051
rect 125823 290023 125851 290051
rect 125637 289961 125665 289989
rect 125699 289961 125727 289989
rect 125761 289961 125789 289989
rect 125823 289961 125851 289989
rect 125637 281147 125665 281175
rect 125699 281147 125727 281175
rect 125761 281147 125789 281175
rect 125823 281147 125851 281175
rect 125637 281085 125665 281113
rect 125699 281085 125727 281113
rect 125761 281085 125789 281113
rect 125823 281085 125851 281113
rect 125637 281023 125665 281051
rect 125699 281023 125727 281051
rect 125761 281023 125789 281051
rect 125823 281023 125851 281051
rect 125637 280961 125665 280989
rect 125699 280961 125727 280989
rect 125761 280961 125789 280989
rect 125823 280961 125851 280989
rect 127497 299058 127525 299086
rect 127559 299058 127587 299086
rect 127621 299058 127649 299086
rect 127683 299058 127711 299086
rect 127497 298996 127525 299024
rect 127559 298996 127587 299024
rect 127621 298996 127649 299024
rect 127683 298996 127711 299024
rect 127497 298934 127525 298962
rect 127559 298934 127587 298962
rect 127621 298934 127649 298962
rect 127683 298934 127711 298962
rect 127497 298872 127525 298900
rect 127559 298872 127587 298900
rect 127621 298872 127649 298900
rect 127683 298872 127711 298900
rect 127497 293147 127525 293175
rect 127559 293147 127587 293175
rect 127621 293147 127649 293175
rect 127683 293147 127711 293175
rect 127497 293085 127525 293113
rect 127559 293085 127587 293113
rect 127621 293085 127649 293113
rect 127683 293085 127711 293113
rect 127497 293023 127525 293051
rect 127559 293023 127587 293051
rect 127621 293023 127649 293051
rect 127683 293023 127711 293051
rect 127497 292961 127525 292989
rect 127559 292961 127587 292989
rect 127621 292961 127649 292989
rect 127683 292961 127711 292989
rect 127497 284147 127525 284175
rect 127559 284147 127587 284175
rect 127621 284147 127649 284175
rect 127683 284147 127711 284175
rect 127497 284085 127525 284113
rect 127559 284085 127587 284113
rect 127621 284085 127649 284113
rect 127683 284085 127711 284113
rect 127497 284023 127525 284051
rect 127559 284023 127587 284051
rect 127621 284023 127649 284051
rect 127683 284023 127711 284051
rect 127497 283961 127525 283989
rect 127559 283961 127587 283989
rect 127621 283961 127649 283989
rect 127683 283961 127711 283989
rect 140997 298578 141025 298606
rect 141059 298578 141087 298606
rect 141121 298578 141149 298606
rect 141183 298578 141211 298606
rect 140997 298516 141025 298544
rect 141059 298516 141087 298544
rect 141121 298516 141149 298544
rect 141183 298516 141211 298544
rect 140997 298454 141025 298482
rect 141059 298454 141087 298482
rect 141121 298454 141149 298482
rect 141183 298454 141211 298482
rect 140997 298392 141025 298420
rect 141059 298392 141087 298420
rect 141121 298392 141149 298420
rect 141183 298392 141211 298420
rect 140997 290147 141025 290175
rect 141059 290147 141087 290175
rect 141121 290147 141149 290175
rect 141183 290147 141211 290175
rect 140997 290085 141025 290113
rect 141059 290085 141087 290113
rect 141121 290085 141149 290113
rect 141183 290085 141211 290113
rect 140997 290023 141025 290051
rect 141059 290023 141087 290051
rect 141121 290023 141149 290051
rect 141183 290023 141211 290051
rect 140997 289961 141025 289989
rect 141059 289961 141087 289989
rect 141121 289961 141149 289989
rect 141183 289961 141211 289989
rect 140997 281147 141025 281175
rect 141059 281147 141087 281175
rect 141121 281147 141149 281175
rect 141183 281147 141211 281175
rect 140997 281085 141025 281113
rect 141059 281085 141087 281113
rect 141121 281085 141149 281113
rect 141183 281085 141211 281113
rect 140997 281023 141025 281051
rect 141059 281023 141087 281051
rect 141121 281023 141149 281051
rect 141183 281023 141211 281051
rect 140997 280961 141025 280989
rect 141059 280961 141087 280989
rect 141121 280961 141149 280989
rect 141183 280961 141211 280989
rect 142857 299058 142885 299086
rect 142919 299058 142947 299086
rect 142981 299058 143009 299086
rect 143043 299058 143071 299086
rect 142857 298996 142885 299024
rect 142919 298996 142947 299024
rect 142981 298996 143009 299024
rect 143043 298996 143071 299024
rect 142857 298934 142885 298962
rect 142919 298934 142947 298962
rect 142981 298934 143009 298962
rect 143043 298934 143071 298962
rect 142857 298872 142885 298900
rect 142919 298872 142947 298900
rect 142981 298872 143009 298900
rect 143043 298872 143071 298900
rect 142857 293147 142885 293175
rect 142919 293147 142947 293175
rect 142981 293147 143009 293175
rect 143043 293147 143071 293175
rect 142857 293085 142885 293113
rect 142919 293085 142947 293113
rect 142981 293085 143009 293113
rect 143043 293085 143071 293113
rect 142857 293023 142885 293051
rect 142919 293023 142947 293051
rect 142981 293023 143009 293051
rect 143043 293023 143071 293051
rect 142857 292961 142885 292989
rect 142919 292961 142947 292989
rect 142981 292961 143009 292989
rect 143043 292961 143071 292989
rect 142857 284147 142885 284175
rect 142919 284147 142947 284175
rect 142981 284147 143009 284175
rect 143043 284147 143071 284175
rect 142857 284085 142885 284113
rect 142919 284085 142947 284113
rect 142981 284085 143009 284113
rect 143043 284085 143071 284113
rect 142857 284023 142885 284051
rect 142919 284023 142947 284051
rect 142981 284023 143009 284051
rect 143043 284023 143071 284051
rect 142857 283961 142885 283989
rect 142919 283961 142947 283989
rect 142981 283961 143009 283989
rect 143043 283961 143071 283989
rect 156357 298578 156385 298606
rect 156419 298578 156447 298606
rect 156481 298578 156509 298606
rect 156543 298578 156571 298606
rect 156357 298516 156385 298544
rect 156419 298516 156447 298544
rect 156481 298516 156509 298544
rect 156543 298516 156571 298544
rect 156357 298454 156385 298482
rect 156419 298454 156447 298482
rect 156481 298454 156509 298482
rect 156543 298454 156571 298482
rect 156357 298392 156385 298420
rect 156419 298392 156447 298420
rect 156481 298392 156509 298420
rect 156543 298392 156571 298420
rect 156357 290147 156385 290175
rect 156419 290147 156447 290175
rect 156481 290147 156509 290175
rect 156543 290147 156571 290175
rect 156357 290085 156385 290113
rect 156419 290085 156447 290113
rect 156481 290085 156509 290113
rect 156543 290085 156571 290113
rect 156357 290023 156385 290051
rect 156419 290023 156447 290051
rect 156481 290023 156509 290051
rect 156543 290023 156571 290051
rect 156357 289961 156385 289989
rect 156419 289961 156447 289989
rect 156481 289961 156509 289989
rect 156543 289961 156571 289989
rect 156357 281147 156385 281175
rect 156419 281147 156447 281175
rect 156481 281147 156509 281175
rect 156543 281147 156571 281175
rect 156357 281085 156385 281113
rect 156419 281085 156447 281113
rect 156481 281085 156509 281113
rect 156543 281085 156571 281113
rect 156357 281023 156385 281051
rect 156419 281023 156447 281051
rect 156481 281023 156509 281051
rect 156543 281023 156571 281051
rect 156357 280961 156385 280989
rect 156419 280961 156447 280989
rect 156481 280961 156509 280989
rect 156543 280961 156571 280989
rect 158217 299058 158245 299086
rect 158279 299058 158307 299086
rect 158341 299058 158369 299086
rect 158403 299058 158431 299086
rect 158217 298996 158245 299024
rect 158279 298996 158307 299024
rect 158341 298996 158369 299024
rect 158403 298996 158431 299024
rect 158217 298934 158245 298962
rect 158279 298934 158307 298962
rect 158341 298934 158369 298962
rect 158403 298934 158431 298962
rect 158217 298872 158245 298900
rect 158279 298872 158307 298900
rect 158341 298872 158369 298900
rect 158403 298872 158431 298900
rect 158217 293147 158245 293175
rect 158279 293147 158307 293175
rect 158341 293147 158369 293175
rect 158403 293147 158431 293175
rect 158217 293085 158245 293113
rect 158279 293085 158307 293113
rect 158341 293085 158369 293113
rect 158403 293085 158431 293113
rect 158217 293023 158245 293051
rect 158279 293023 158307 293051
rect 158341 293023 158369 293051
rect 158403 293023 158431 293051
rect 158217 292961 158245 292989
rect 158279 292961 158307 292989
rect 158341 292961 158369 292989
rect 158403 292961 158431 292989
rect 158217 284147 158245 284175
rect 158279 284147 158307 284175
rect 158341 284147 158369 284175
rect 158403 284147 158431 284175
rect 158217 284085 158245 284113
rect 158279 284085 158307 284113
rect 158341 284085 158369 284113
rect 158403 284085 158431 284113
rect 158217 284023 158245 284051
rect 158279 284023 158307 284051
rect 158341 284023 158369 284051
rect 158403 284023 158431 284051
rect 158217 283961 158245 283989
rect 158279 283961 158307 283989
rect 158341 283961 158369 283989
rect 158403 283961 158431 283989
rect 171717 298578 171745 298606
rect 171779 298578 171807 298606
rect 171841 298578 171869 298606
rect 171903 298578 171931 298606
rect 171717 298516 171745 298544
rect 171779 298516 171807 298544
rect 171841 298516 171869 298544
rect 171903 298516 171931 298544
rect 171717 298454 171745 298482
rect 171779 298454 171807 298482
rect 171841 298454 171869 298482
rect 171903 298454 171931 298482
rect 171717 298392 171745 298420
rect 171779 298392 171807 298420
rect 171841 298392 171869 298420
rect 171903 298392 171931 298420
rect 171717 290147 171745 290175
rect 171779 290147 171807 290175
rect 171841 290147 171869 290175
rect 171903 290147 171931 290175
rect 171717 290085 171745 290113
rect 171779 290085 171807 290113
rect 171841 290085 171869 290113
rect 171903 290085 171931 290113
rect 171717 290023 171745 290051
rect 171779 290023 171807 290051
rect 171841 290023 171869 290051
rect 171903 290023 171931 290051
rect 171717 289961 171745 289989
rect 171779 289961 171807 289989
rect 171841 289961 171869 289989
rect 171903 289961 171931 289989
rect 171717 281147 171745 281175
rect 171779 281147 171807 281175
rect 171841 281147 171869 281175
rect 171903 281147 171931 281175
rect 171717 281085 171745 281113
rect 171779 281085 171807 281113
rect 171841 281085 171869 281113
rect 171903 281085 171931 281113
rect 171717 281023 171745 281051
rect 171779 281023 171807 281051
rect 171841 281023 171869 281051
rect 171903 281023 171931 281051
rect 171717 280961 171745 280989
rect 171779 280961 171807 280989
rect 171841 280961 171869 280989
rect 171903 280961 171931 280989
rect 173577 299058 173605 299086
rect 173639 299058 173667 299086
rect 173701 299058 173729 299086
rect 173763 299058 173791 299086
rect 173577 298996 173605 299024
rect 173639 298996 173667 299024
rect 173701 298996 173729 299024
rect 173763 298996 173791 299024
rect 173577 298934 173605 298962
rect 173639 298934 173667 298962
rect 173701 298934 173729 298962
rect 173763 298934 173791 298962
rect 173577 298872 173605 298900
rect 173639 298872 173667 298900
rect 173701 298872 173729 298900
rect 173763 298872 173791 298900
rect 173577 293147 173605 293175
rect 173639 293147 173667 293175
rect 173701 293147 173729 293175
rect 173763 293147 173791 293175
rect 173577 293085 173605 293113
rect 173639 293085 173667 293113
rect 173701 293085 173729 293113
rect 173763 293085 173791 293113
rect 173577 293023 173605 293051
rect 173639 293023 173667 293051
rect 173701 293023 173729 293051
rect 173763 293023 173791 293051
rect 173577 292961 173605 292989
rect 173639 292961 173667 292989
rect 173701 292961 173729 292989
rect 173763 292961 173791 292989
rect 173577 284147 173605 284175
rect 173639 284147 173667 284175
rect 173701 284147 173729 284175
rect 173763 284147 173791 284175
rect 173577 284085 173605 284113
rect 173639 284085 173667 284113
rect 173701 284085 173729 284113
rect 173763 284085 173791 284113
rect 173577 284023 173605 284051
rect 173639 284023 173667 284051
rect 173701 284023 173729 284051
rect 173763 284023 173791 284051
rect 173577 283961 173605 283989
rect 173639 283961 173667 283989
rect 173701 283961 173729 283989
rect 173763 283961 173791 283989
rect 187077 298578 187105 298606
rect 187139 298578 187167 298606
rect 187201 298578 187229 298606
rect 187263 298578 187291 298606
rect 187077 298516 187105 298544
rect 187139 298516 187167 298544
rect 187201 298516 187229 298544
rect 187263 298516 187291 298544
rect 187077 298454 187105 298482
rect 187139 298454 187167 298482
rect 187201 298454 187229 298482
rect 187263 298454 187291 298482
rect 187077 298392 187105 298420
rect 187139 298392 187167 298420
rect 187201 298392 187229 298420
rect 187263 298392 187291 298420
rect 187077 290147 187105 290175
rect 187139 290147 187167 290175
rect 187201 290147 187229 290175
rect 187263 290147 187291 290175
rect 187077 290085 187105 290113
rect 187139 290085 187167 290113
rect 187201 290085 187229 290113
rect 187263 290085 187291 290113
rect 187077 290023 187105 290051
rect 187139 290023 187167 290051
rect 187201 290023 187229 290051
rect 187263 290023 187291 290051
rect 187077 289961 187105 289989
rect 187139 289961 187167 289989
rect 187201 289961 187229 289989
rect 187263 289961 187291 289989
rect 187077 281147 187105 281175
rect 187139 281147 187167 281175
rect 187201 281147 187229 281175
rect 187263 281147 187291 281175
rect 187077 281085 187105 281113
rect 187139 281085 187167 281113
rect 187201 281085 187229 281113
rect 187263 281085 187291 281113
rect 187077 281023 187105 281051
rect 187139 281023 187167 281051
rect 187201 281023 187229 281051
rect 187263 281023 187291 281051
rect 187077 280961 187105 280989
rect 187139 280961 187167 280989
rect 187201 280961 187229 280989
rect 187263 280961 187291 280989
rect 188937 299058 188965 299086
rect 188999 299058 189027 299086
rect 189061 299058 189089 299086
rect 189123 299058 189151 299086
rect 188937 298996 188965 299024
rect 188999 298996 189027 299024
rect 189061 298996 189089 299024
rect 189123 298996 189151 299024
rect 188937 298934 188965 298962
rect 188999 298934 189027 298962
rect 189061 298934 189089 298962
rect 189123 298934 189151 298962
rect 188937 298872 188965 298900
rect 188999 298872 189027 298900
rect 189061 298872 189089 298900
rect 189123 298872 189151 298900
rect 188937 293147 188965 293175
rect 188999 293147 189027 293175
rect 189061 293147 189089 293175
rect 189123 293147 189151 293175
rect 188937 293085 188965 293113
rect 188999 293085 189027 293113
rect 189061 293085 189089 293113
rect 189123 293085 189151 293113
rect 188937 293023 188965 293051
rect 188999 293023 189027 293051
rect 189061 293023 189089 293051
rect 189123 293023 189151 293051
rect 188937 292961 188965 292989
rect 188999 292961 189027 292989
rect 189061 292961 189089 292989
rect 189123 292961 189151 292989
rect 188937 284147 188965 284175
rect 188999 284147 189027 284175
rect 189061 284147 189089 284175
rect 189123 284147 189151 284175
rect 188937 284085 188965 284113
rect 188999 284085 189027 284113
rect 189061 284085 189089 284113
rect 189123 284085 189151 284113
rect 188937 284023 188965 284051
rect 188999 284023 189027 284051
rect 189061 284023 189089 284051
rect 189123 284023 189151 284051
rect 188937 283961 188965 283989
rect 188999 283961 189027 283989
rect 189061 283961 189089 283989
rect 189123 283961 189151 283989
rect 202437 298578 202465 298606
rect 202499 298578 202527 298606
rect 202561 298578 202589 298606
rect 202623 298578 202651 298606
rect 202437 298516 202465 298544
rect 202499 298516 202527 298544
rect 202561 298516 202589 298544
rect 202623 298516 202651 298544
rect 202437 298454 202465 298482
rect 202499 298454 202527 298482
rect 202561 298454 202589 298482
rect 202623 298454 202651 298482
rect 202437 298392 202465 298420
rect 202499 298392 202527 298420
rect 202561 298392 202589 298420
rect 202623 298392 202651 298420
rect 202437 290147 202465 290175
rect 202499 290147 202527 290175
rect 202561 290147 202589 290175
rect 202623 290147 202651 290175
rect 202437 290085 202465 290113
rect 202499 290085 202527 290113
rect 202561 290085 202589 290113
rect 202623 290085 202651 290113
rect 202437 290023 202465 290051
rect 202499 290023 202527 290051
rect 202561 290023 202589 290051
rect 202623 290023 202651 290051
rect 202437 289961 202465 289989
rect 202499 289961 202527 289989
rect 202561 289961 202589 289989
rect 202623 289961 202651 289989
rect 202437 281147 202465 281175
rect 202499 281147 202527 281175
rect 202561 281147 202589 281175
rect 202623 281147 202651 281175
rect 202437 281085 202465 281113
rect 202499 281085 202527 281113
rect 202561 281085 202589 281113
rect 202623 281085 202651 281113
rect 202437 281023 202465 281051
rect 202499 281023 202527 281051
rect 202561 281023 202589 281051
rect 202623 281023 202651 281051
rect 202437 280961 202465 280989
rect 202499 280961 202527 280989
rect 202561 280961 202589 280989
rect 202623 280961 202651 280989
rect 204297 299058 204325 299086
rect 204359 299058 204387 299086
rect 204421 299058 204449 299086
rect 204483 299058 204511 299086
rect 204297 298996 204325 299024
rect 204359 298996 204387 299024
rect 204421 298996 204449 299024
rect 204483 298996 204511 299024
rect 204297 298934 204325 298962
rect 204359 298934 204387 298962
rect 204421 298934 204449 298962
rect 204483 298934 204511 298962
rect 204297 298872 204325 298900
rect 204359 298872 204387 298900
rect 204421 298872 204449 298900
rect 204483 298872 204511 298900
rect 204297 293147 204325 293175
rect 204359 293147 204387 293175
rect 204421 293147 204449 293175
rect 204483 293147 204511 293175
rect 204297 293085 204325 293113
rect 204359 293085 204387 293113
rect 204421 293085 204449 293113
rect 204483 293085 204511 293113
rect 204297 293023 204325 293051
rect 204359 293023 204387 293051
rect 204421 293023 204449 293051
rect 204483 293023 204511 293051
rect 204297 292961 204325 292989
rect 204359 292961 204387 292989
rect 204421 292961 204449 292989
rect 204483 292961 204511 292989
rect 204297 284147 204325 284175
rect 204359 284147 204387 284175
rect 204421 284147 204449 284175
rect 204483 284147 204511 284175
rect 204297 284085 204325 284113
rect 204359 284085 204387 284113
rect 204421 284085 204449 284113
rect 204483 284085 204511 284113
rect 204297 284023 204325 284051
rect 204359 284023 204387 284051
rect 204421 284023 204449 284051
rect 204483 284023 204511 284051
rect 204297 283961 204325 283989
rect 204359 283961 204387 283989
rect 204421 283961 204449 283989
rect 204483 283961 204511 283989
rect 217797 298578 217825 298606
rect 217859 298578 217887 298606
rect 217921 298578 217949 298606
rect 217983 298578 218011 298606
rect 217797 298516 217825 298544
rect 217859 298516 217887 298544
rect 217921 298516 217949 298544
rect 217983 298516 218011 298544
rect 217797 298454 217825 298482
rect 217859 298454 217887 298482
rect 217921 298454 217949 298482
rect 217983 298454 218011 298482
rect 217797 298392 217825 298420
rect 217859 298392 217887 298420
rect 217921 298392 217949 298420
rect 217983 298392 218011 298420
rect 217797 290147 217825 290175
rect 217859 290147 217887 290175
rect 217921 290147 217949 290175
rect 217983 290147 218011 290175
rect 217797 290085 217825 290113
rect 217859 290085 217887 290113
rect 217921 290085 217949 290113
rect 217983 290085 218011 290113
rect 217797 290023 217825 290051
rect 217859 290023 217887 290051
rect 217921 290023 217949 290051
rect 217983 290023 218011 290051
rect 217797 289961 217825 289989
rect 217859 289961 217887 289989
rect 217921 289961 217949 289989
rect 217983 289961 218011 289989
rect 217797 281147 217825 281175
rect 217859 281147 217887 281175
rect 217921 281147 217949 281175
rect 217983 281147 218011 281175
rect 217797 281085 217825 281113
rect 217859 281085 217887 281113
rect 217921 281085 217949 281113
rect 217983 281085 218011 281113
rect 217797 281023 217825 281051
rect 217859 281023 217887 281051
rect 217921 281023 217949 281051
rect 217983 281023 218011 281051
rect 217797 280961 217825 280989
rect 217859 280961 217887 280989
rect 217921 280961 217949 280989
rect 217983 280961 218011 280989
rect 219657 299058 219685 299086
rect 219719 299058 219747 299086
rect 219781 299058 219809 299086
rect 219843 299058 219871 299086
rect 219657 298996 219685 299024
rect 219719 298996 219747 299024
rect 219781 298996 219809 299024
rect 219843 298996 219871 299024
rect 219657 298934 219685 298962
rect 219719 298934 219747 298962
rect 219781 298934 219809 298962
rect 219843 298934 219871 298962
rect 219657 298872 219685 298900
rect 219719 298872 219747 298900
rect 219781 298872 219809 298900
rect 219843 298872 219871 298900
rect 219657 293147 219685 293175
rect 219719 293147 219747 293175
rect 219781 293147 219809 293175
rect 219843 293147 219871 293175
rect 219657 293085 219685 293113
rect 219719 293085 219747 293113
rect 219781 293085 219809 293113
rect 219843 293085 219871 293113
rect 219657 293023 219685 293051
rect 219719 293023 219747 293051
rect 219781 293023 219809 293051
rect 219843 293023 219871 293051
rect 219657 292961 219685 292989
rect 219719 292961 219747 292989
rect 219781 292961 219809 292989
rect 219843 292961 219871 292989
rect 219657 284147 219685 284175
rect 219719 284147 219747 284175
rect 219781 284147 219809 284175
rect 219843 284147 219871 284175
rect 219657 284085 219685 284113
rect 219719 284085 219747 284113
rect 219781 284085 219809 284113
rect 219843 284085 219871 284113
rect 219657 284023 219685 284051
rect 219719 284023 219747 284051
rect 219781 284023 219809 284051
rect 219843 284023 219871 284051
rect 219657 283961 219685 283989
rect 219719 283961 219747 283989
rect 219781 283961 219809 283989
rect 219843 283961 219871 283989
rect 233157 298578 233185 298606
rect 233219 298578 233247 298606
rect 233281 298578 233309 298606
rect 233343 298578 233371 298606
rect 233157 298516 233185 298544
rect 233219 298516 233247 298544
rect 233281 298516 233309 298544
rect 233343 298516 233371 298544
rect 233157 298454 233185 298482
rect 233219 298454 233247 298482
rect 233281 298454 233309 298482
rect 233343 298454 233371 298482
rect 233157 298392 233185 298420
rect 233219 298392 233247 298420
rect 233281 298392 233309 298420
rect 233343 298392 233371 298420
rect 233157 290147 233185 290175
rect 233219 290147 233247 290175
rect 233281 290147 233309 290175
rect 233343 290147 233371 290175
rect 233157 290085 233185 290113
rect 233219 290085 233247 290113
rect 233281 290085 233309 290113
rect 233343 290085 233371 290113
rect 233157 290023 233185 290051
rect 233219 290023 233247 290051
rect 233281 290023 233309 290051
rect 233343 290023 233371 290051
rect 233157 289961 233185 289989
rect 233219 289961 233247 289989
rect 233281 289961 233309 289989
rect 233343 289961 233371 289989
rect 233157 281147 233185 281175
rect 233219 281147 233247 281175
rect 233281 281147 233309 281175
rect 233343 281147 233371 281175
rect 233157 281085 233185 281113
rect 233219 281085 233247 281113
rect 233281 281085 233309 281113
rect 233343 281085 233371 281113
rect 233157 281023 233185 281051
rect 233219 281023 233247 281051
rect 233281 281023 233309 281051
rect 233343 281023 233371 281051
rect 233157 280961 233185 280989
rect 233219 280961 233247 280989
rect 233281 280961 233309 280989
rect 233343 280961 233371 280989
rect 235017 299058 235045 299086
rect 235079 299058 235107 299086
rect 235141 299058 235169 299086
rect 235203 299058 235231 299086
rect 235017 298996 235045 299024
rect 235079 298996 235107 299024
rect 235141 298996 235169 299024
rect 235203 298996 235231 299024
rect 235017 298934 235045 298962
rect 235079 298934 235107 298962
rect 235141 298934 235169 298962
rect 235203 298934 235231 298962
rect 235017 298872 235045 298900
rect 235079 298872 235107 298900
rect 235141 298872 235169 298900
rect 235203 298872 235231 298900
rect 235017 293147 235045 293175
rect 235079 293147 235107 293175
rect 235141 293147 235169 293175
rect 235203 293147 235231 293175
rect 235017 293085 235045 293113
rect 235079 293085 235107 293113
rect 235141 293085 235169 293113
rect 235203 293085 235231 293113
rect 235017 293023 235045 293051
rect 235079 293023 235107 293051
rect 235141 293023 235169 293051
rect 235203 293023 235231 293051
rect 235017 292961 235045 292989
rect 235079 292961 235107 292989
rect 235141 292961 235169 292989
rect 235203 292961 235231 292989
rect 235017 284147 235045 284175
rect 235079 284147 235107 284175
rect 235141 284147 235169 284175
rect 235203 284147 235231 284175
rect 235017 284085 235045 284113
rect 235079 284085 235107 284113
rect 235141 284085 235169 284113
rect 235203 284085 235231 284113
rect 235017 284023 235045 284051
rect 235079 284023 235107 284051
rect 235141 284023 235169 284051
rect 235203 284023 235231 284051
rect 235017 283961 235045 283989
rect 235079 283961 235107 283989
rect 235141 283961 235169 283989
rect 235203 283961 235231 283989
rect 248517 298578 248545 298606
rect 248579 298578 248607 298606
rect 248641 298578 248669 298606
rect 248703 298578 248731 298606
rect 248517 298516 248545 298544
rect 248579 298516 248607 298544
rect 248641 298516 248669 298544
rect 248703 298516 248731 298544
rect 248517 298454 248545 298482
rect 248579 298454 248607 298482
rect 248641 298454 248669 298482
rect 248703 298454 248731 298482
rect 248517 298392 248545 298420
rect 248579 298392 248607 298420
rect 248641 298392 248669 298420
rect 248703 298392 248731 298420
rect 248517 290147 248545 290175
rect 248579 290147 248607 290175
rect 248641 290147 248669 290175
rect 248703 290147 248731 290175
rect 248517 290085 248545 290113
rect 248579 290085 248607 290113
rect 248641 290085 248669 290113
rect 248703 290085 248731 290113
rect 248517 290023 248545 290051
rect 248579 290023 248607 290051
rect 248641 290023 248669 290051
rect 248703 290023 248731 290051
rect 248517 289961 248545 289989
rect 248579 289961 248607 289989
rect 248641 289961 248669 289989
rect 248703 289961 248731 289989
rect 248517 281147 248545 281175
rect 248579 281147 248607 281175
rect 248641 281147 248669 281175
rect 248703 281147 248731 281175
rect 248517 281085 248545 281113
rect 248579 281085 248607 281113
rect 248641 281085 248669 281113
rect 248703 281085 248731 281113
rect 248517 281023 248545 281051
rect 248579 281023 248607 281051
rect 248641 281023 248669 281051
rect 248703 281023 248731 281051
rect 248517 280961 248545 280989
rect 248579 280961 248607 280989
rect 248641 280961 248669 280989
rect 248703 280961 248731 280989
rect 250377 299058 250405 299086
rect 250439 299058 250467 299086
rect 250501 299058 250529 299086
rect 250563 299058 250591 299086
rect 250377 298996 250405 299024
rect 250439 298996 250467 299024
rect 250501 298996 250529 299024
rect 250563 298996 250591 299024
rect 250377 298934 250405 298962
rect 250439 298934 250467 298962
rect 250501 298934 250529 298962
rect 250563 298934 250591 298962
rect 250377 298872 250405 298900
rect 250439 298872 250467 298900
rect 250501 298872 250529 298900
rect 250563 298872 250591 298900
rect 250377 293147 250405 293175
rect 250439 293147 250467 293175
rect 250501 293147 250529 293175
rect 250563 293147 250591 293175
rect 250377 293085 250405 293113
rect 250439 293085 250467 293113
rect 250501 293085 250529 293113
rect 250563 293085 250591 293113
rect 250377 293023 250405 293051
rect 250439 293023 250467 293051
rect 250501 293023 250529 293051
rect 250563 293023 250591 293051
rect 250377 292961 250405 292989
rect 250439 292961 250467 292989
rect 250501 292961 250529 292989
rect 250563 292961 250591 292989
rect 250377 284147 250405 284175
rect 250439 284147 250467 284175
rect 250501 284147 250529 284175
rect 250563 284147 250591 284175
rect 250377 284085 250405 284113
rect 250439 284085 250467 284113
rect 250501 284085 250529 284113
rect 250563 284085 250591 284113
rect 250377 284023 250405 284051
rect 250439 284023 250467 284051
rect 250501 284023 250529 284051
rect 250563 284023 250591 284051
rect 250377 283961 250405 283989
rect 250439 283961 250467 283989
rect 250501 283961 250529 283989
rect 250563 283961 250591 283989
rect 263877 298578 263905 298606
rect 263939 298578 263967 298606
rect 264001 298578 264029 298606
rect 264063 298578 264091 298606
rect 263877 298516 263905 298544
rect 263939 298516 263967 298544
rect 264001 298516 264029 298544
rect 264063 298516 264091 298544
rect 263877 298454 263905 298482
rect 263939 298454 263967 298482
rect 264001 298454 264029 298482
rect 264063 298454 264091 298482
rect 263877 298392 263905 298420
rect 263939 298392 263967 298420
rect 264001 298392 264029 298420
rect 264063 298392 264091 298420
rect 263877 290147 263905 290175
rect 263939 290147 263967 290175
rect 264001 290147 264029 290175
rect 264063 290147 264091 290175
rect 263877 290085 263905 290113
rect 263939 290085 263967 290113
rect 264001 290085 264029 290113
rect 264063 290085 264091 290113
rect 263877 290023 263905 290051
rect 263939 290023 263967 290051
rect 264001 290023 264029 290051
rect 264063 290023 264091 290051
rect 263877 289961 263905 289989
rect 263939 289961 263967 289989
rect 264001 289961 264029 289989
rect 264063 289961 264091 289989
rect 263877 281147 263905 281175
rect 263939 281147 263967 281175
rect 264001 281147 264029 281175
rect 264063 281147 264091 281175
rect 263877 281085 263905 281113
rect 263939 281085 263967 281113
rect 264001 281085 264029 281113
rect 264063 281085 264091 281113
rect 263877 281023 263905 281051
rect 263939 281023 263967 281051
rect 264001 281023 264029 281051
rect 264063 281023 264091 281051
rect 263877 280961 263905 280989
rect 263939 280961 263967 280989
rect 264001 280961 264029 280989
rect 264063 280961 264091 280989
rect 265737 299058 265765 299086
rect 265799 299058 265827 299086
rect 265861 299058 265889 299086
rect 265923 299058 265951 299086
rect 265737 298996 265765 299024
rect 265799 298996 265827 299024
rect 265861 298996 265889 299024
rect 265923 298996 265951 299024
rect 265737 298934 265765 298962
rect 265799 298934 265827 298962
rect 265861 298934 265889 298962
rect 265923 298934 265951 298962
rect 265737 298872 265765 298900
rect 265799 298872 265827 298900
rect 265861 298872 265889 298900
rect 265923 298872 265951 298900
rect 265737 293147 265765 293175
rect 265799 293147 265827 293175
rect 265861 293147 265889 293175
rect 265923 293147 265951 293175
rect 265737 293085 265765 293113
rect 265799 293085 265827 293113
rect 265861 293085 265889 293113
rect 265923 293085 265951 293113
rect 265737 293023 265765 293051
rect 265799 293023 265827 293051
rect 265861 293023 265889 293051
rect 265923 293023 265951 293051
rect 265737 292961 265765 292989
rect 265799 292961 265827 292989
rect 265861 292961 265889 292989
rect 265923 292961 265951 292989
rect 265737 284147 265765 284175
rect 265799 284147 265827 284175
rect 265861 284147 265889 284175
rect 265923 284147 265951 284175
rect 265737 284085 265765 284113
rect 265799 284085 265827 284113
rect 265861 284085 265889 284113
rect 265923 284085 265951 284113
rect 265737 284023 265765 284051
rect 265799 284023 265827 284051
rect 265861 284023 265889 284051
rect 265923 284023 265951 284051
rect 265737 283961 265765 283989
rect 265799 283961 265827 283989
rect 265861 283961 265889 283989
rect 265923 283961 265951 283989
rect 279237 298578 279265 298606
rect 279299 298578 279327 298606
rect 279361 298578 279389 298606
rect 279423 298578 279451 298606
rect 279237 298516 279265 298544
rect 279299 298516 279327 298544
rect 279361 298516 279389 298544
rect 279423 298516 279451 298544
rect 279237 298454 279265 298482
rect 279299 298454 279327 298482
rect 279361 298454 279389 298482
rect 279423 298454 279451 298482
rect 279237 298392 279265 298420
rect 279299 298392 279327 298420
rect 279361 298392 279389 298420
rect 279423 298392 279451 298420
rect 279237 290147 279265 290175
rect 279299 290147 279327 290175
rect 279361 290147 279389 290175
rect 279423 290147 279451 290175
rect 279237 290085 279265 290113
rect 279299 290085 279327 290113
rect 279361 290085 279389 290113
rect 279423 290085 279451 290113
rect 279237 290023 279265 290051
rect 279299 290023 279327 290051
rect 279361 290023 279389 290051
rect 279423 290023 279451 290051
rect 279237 289961 279265 289989
rect 279299 289961 279327 289989
rect 279361 289961 279389 289989
rect 279423 289961 279451 289989
rect 279237 281147 279265 281175
rect 279299 281147 279327 281175
rect 279361 281147 279389 281175
rect 279423 281147 279451 281175
rect 279237 281085 279265 281113
rect 279299 281085 279327 281113
rect 279361 281085 279389 281113
rect 279423 281085 279451 281113
rect 279237 281023 279265 281051
rect 279299 281023 279327 281051
rect 279361 281023 279389 281051
rect 279423 281023 279451 281051
rect 279237 280961 279265 280989
rect 279299 280961 279327 280989
rect 279361 280961 279389 280989
rect 279423 280961 279451 280989
rect 96777 275147 96805 275175
rect 96839 275147 96867 275175
rect 96901 275147 96929 275175
rect 96963 275147 96991 275175
rect 96777 275085 96805 275113
rect 96839 275085 96867 275113
rect 96901 275085 96929 275113
rect 96963 275085 96991 275113
rect 96777 275023 96805 275051
rect 96839 275023 96867 275051
rect 96901 275023 96929 275051
rect 96963 275023 96991 275051
rect 109939 275147 109967 275175
rect 110001 275147 110029 275175
rect 109939 275085 109967 275113
rect 110001 275085 110029 275113
rect 109939 275023 109967 275051
rect 110001 275023 110029 275051
rect 96777 274961 96805 274989
rect 96839 274961 96867 274989
rect 96901 274961 96929 274989
rect 96963 274961 96991 274989
rect 96777 266147 96805 266175
rect 96839 266147 96867 266175
rect 96901 266147 96929 266175
rect 96963 266147 96991 266175
rect 96777 266085 96805 266113
rect 96839 266085 96867 266113
rect 96901 266085 96929 266113
rect 96963 266085 96991 266113
rect 96777 266023 96805 266051
rect 96839 266023 96867 266051
rect 96901 266023 96929 266051
rect 96963 266023 96991 266051
rect 96777 265961 96805 265989
rect 96839 265961 96867 265989
rect 96901 265961 96929 265989
rect 96963 265961 96991 265989
rect 96777 257147 96805 257175
rect 96839 257147 96867 257175
rect 96901 257147 96929 257175
rect 96963 257147 96991 257175
rect 96777 257085 96805 257113
rect 96839 257085 96867 257113
rect 96901 257085 96929 257113
rect 96963 257085 96991 257113
rect 96777 257023 96805 257051
rect 96839 257023 96867 257051
rect 96901 257023 96929 257051
rect 96963 257023 96991 257051
rect 96777 256961 96805 256989
rect 96839 256961 96867 256989
rect 96901 256961 96929 256989
rect 96963 256961 96991 256989
rect 96777 248147 96805 248175
rect 96839 248147 96867 248175
rect 96901 248147 96929 248175
rect 96963 248147 96991 248175
rect 96777 248085 96805 248113
rect 96839 248085 96867 248113
rect 96901 248085 96929 248113
rect 96963 248085 96991 248113
rect 96777 248023 96805 248051
rect 96839 248023 96867 248051
rect 96901 248023 96929 248051
rect 96963 248023 96991 248051
rect 96777 247961 96805 247989
rect 96839 247961 96867 247989
rect 96901 247961 96929 247989
rect 96963 247961 96991 247989
rect 96777 239147 96805 239175
rect 96839 239147 96867 239175
rect 96901 239147 96929 239175
rect 96963 239147 96991 239175
rect 96777 239085 96805 239113
rect 96839 239085 96867 239113
rect 96901 239085 96929 239113
rect 96963 239085 96991 239113
rect 96777 239023 96805 239051
rect 96839 239023 96867 239051
rect 96901 239023 96929 239051
rect 96963 239023 96991 239051
rect 96777 238961 96805 238989
rect 96839 238961 96867 238989
rect 96901 238961 96929 238989
rect 96963 238961 96991 238989
rect 96777 230147 96805 230175
rect 96839 230147 96867 230175
rect 96901 230147 96929 230175
rect 96963 230147 96991 230175
rect 96777 230085 96805 230113
rect 96839 230085 96867 230113
rect 96901 230085 96929 230113
rect 96963 230085 96991 230113
rect 96777 230023 96805 230051
rect 96839 230023 96867 230051
rect 96901 230023 96929 230051
rect 96963 230023 96991 230051
rect 96777 229961 96805 229989
rect 96839 229961 96867 229989
rect 96901 229961 96929 229989
rect 96963 229961 96991 229989
rect 96777 221147 96805 221175
rect 96839 221147 96867 221175
rect 96901 221147 96929 221175
rect 96963 221147 96991 221175
rect 96777 221085 96805 221113
rect 96839 221085 96867 221113
rect 96901 221085 96929 221113
rect 96963 221085 96991 221113
rect 96777 221023 96805 221051
rect 96839 221023 96867 221051
rect 96901 221023 96929 221051
rect 96963 221023 96991 221051
rect 96777 220961 96805 220989
rect 96839 220961 96867 220989
rect 96901 220961 96929 220989
rect 96963 220961 96991 220989
rect 96777 212147 96805 212175
rect 96839 212147 96867 212175
rect 96901 212147 96929 212175
rect 96963 212147 96991 212175
rect 96777 212085 96805 212113
rect 96839 212085 96867 212113
rect 96901 212085 96929 212113
rect 96963 212085 96991 212113
rect 96777 212023 96805 212051
rect 96839 212023 96867 212051
rect 96901 212023 96929 212051
rect 96963 212023 96991 212051
rect 96777 211961 96805 211989
rect 96839 211961 96867 211989
rect 96901 211961 96929 211989
rect 96963 211961 96991 211989
rect 96777 203147 96805 203175
rect 96839 203147 96867 203175
rect 96901 203147 96929 203175
rect 96963 203147 96991 203175
rect 96777 203085 96805 203113
rect 96839 203085 96867 203113
rect 96901 203085 96929 203113
rect 96963 203085 96991 203113
rect 96777 203023 96805 203051
rect 96839 203023 96867 203051
rect 96901 203023 96929 203051
rect 96963 203023 96991 203051
rect 96777 202961 96805 202989
rect 96839 202961 96867 202989
rect 96901 202961 96929 202989
rect 96963 202961 96991 202989
rect 96777 194147 96805 194175
rect 96839 194147 96867 194175
rect 96901 194147 96929 194175
rect 96963 194147 96991 194175
rect 96777 194085 96805 194113
rect 96839 194085 96867 194113
rect 96901 194085 96929 194113
rect 96963 194085 96991 194113
rect 96777 194023 96805 194051
rect 96839 194023 96867 194051
rect 96901 194023 96929 194051
rect 96963 194023 96991 194051
rect 96777 193961 96805 193989
rect 96839 193961 96867 193989
rect 96901 193961 96929 193989
rect 96963 193961 96991 193989
rect 96777 185147 96805 185175
rect 96839 185147 96867 185175
rect 96901 185147 96929 185175
rect 96963 185147 96991 185175
rect 96777 185085 96805 185113
rect 96839 185085 96867 185113
rect 96901 185085 96929 185113
rect 96963 185085 96991 185113
rect 96777 185023 96805 185051
rect 96839 185023 96867 185051
rect 96901 185023 96929 185051
rect 96963 185023 96991 185051
rect 96777 184961 96805 184989
rect 96839 184961 96867 184989
rect 96901 184961 96929 184989
rect 96963 184961 96991 184989
rect 96777 176147 96805 176175
rect 96839 176147 96867 176175
rect 96901 176147 96929 176175
rect 96963 176147 96991 176175
rect 96777 176085 96805 176113
rect 96839 176085 96867 176113
rect 96901 176085 96929 176113
rect 96963 176085 96991 176113
rect 96777 176023 96805 176051
rect 96839 176023 96867 176051
rect 96901 176023 96929 176051
rect 96963 176023 96991 176051
rect 96777 175961 96805 175989
rect 96839 175961 96867 175989
rect 96901 175961 96929 175989
rect 96963 175961 96991 175989
rect 96777 167147 96805 167175
rect 96839 167147 96867 167175
rect 96901 167147 96929 167175
rect 96963 167147 96991 167175
rect 96777 167085 96805 167113
rect 96839 167085 96867 167113
rect 96901 167085 96929 167113
rect 96963 167085 96991 167113
rect 96777 167023 96805 167051
rect 96839 167023 96867 167051
rect 96901 167023 96929 167051
rect 96963 167023 96991 167051
rect 96777 166961 96805 166989
rect 96839 166961 96867 166989
rect 96901 166961 96929 166989
rect 96963 166961 96991 166989
rect 96777 158147 96805 158175
rect 96839 158147 96867 158175
rect 96901 158147 96929 158175
rect 96963 158147 96991 158175
rect 96777 158085 96805 158113
rect 96839 158085 96867 158113
rect 96901 158085 96929 158113
rect 96963 158085 96991 158113
rect 96777 158023 96805 158051
rect 96839 158023 96867 158051
rect 96901 158023 96929 158051
rect 96963 158023 96991 158051
rect 96777 157961 96805 157989
rect 96839 157961 96867 157989
rect 96901 157961 96929 157989
rect 96963 157961 96991 157989
rect 96777 149147 96805 149175
rect 96839 149147 96867 149175
rect 96901 149147 96929 149175
rect 96963 149147 96991 149175
rect 96777 149085 96805 149113
rect 96839 149085 96867 149113
rect 96901 149085 96929 149113
rect 96963 149085 96991 149113
rect 96777 149023 96805 149051
rect 96839 149023 96867 149051
rect 96901 149023 96929 149051
rect 96963 149023 96991 149051
rect 96777 148961 96805 148989
rect 96839 148961 96867 148989
rect 96901 148961 96929 148989
rect 96963 148961 96991 148989
rect 96777 140147 96805 140175
rect 96839 140147 96867 140175
rect 96901 140147 96929 140175
rect 96963 140147 96991 140175
rect 96777 140085 96805 140113
rect 96839 140085 96867 140113
rect 96901 140085 96929 140113
rect 96963 140085 96991 140113
rect 96777 140023 96805 140051
rect 96839 140023 96867 140051
rect 96901 140023 96929 140051
rect 96963 140023 96991 140051
rect 96777 139961 96805 139989
rect 96839 139961 96867 139989
rect 96901 139961 96929 139989
rect 96963 139961 96991 139989
rect 96777 131147 96805 131175
rect 96839 131147 96867 131175
rect 96901 131147 96929 131175
rect 96963 131147 96991 131175
rect 96777 131085 96805 131113
rect 96839 131085 96867 131113
rect 96901 131085 96929 131113
rect 96963 131085 96991 131113
rect 96777 131023 96805 131051
rect 96839 131023 96867 131051
rect 96901 131023 96929 131051
rect 96963 131023 96991 131051
rect 96777 130961 96805 130989
rect 96839 130961 96867 130989
rect 96901 130961 96929 130989
rect 96963 130961 96991 130989
rect 96777 122147 96805 122175
rect 96839 122147 96867 122175
rect 96901 122147 96929 122175
rect 96963 122147 96991 122175
rect 96777 122085 96805 122113
rect 96839 122085 96867 122113
rect 96901 122085 96929 122113
rect 96963 122085 96991 122113
rect 96777 122023 96805 122051
rect 96839 122023 96867 122051
rect 96901 122023 96929 122051
rect 96963 122023 96991 122051
rect 96777 121961 96805 121989
rect 96839 121961 96867 121989
rect 96901 121961 96929 121989
rect 96963 121961 96991 121989
rect 96777 113147 96805 113175
rect 96839 113147 96867 113175
rect 96901 113147 96929 113175
rect 96963 113147 96991 113175
rect 96777 113085 96805 113113
rect 96839 113085 96867 113113
rect 96901 113085 96929 113113
rect 96963 113085 96991 113113
rect 96777 113023 96805 113051
rect 96839 113023 96867 113051
rect 96901 113023 96929 113051
rect 96963 113023 96991 113051
rect 96777 112961 96805 112989
rect 96839 112961 96867 112989
rect 96901 112961 96929 112989
rect 96963 112961 96991 112989
rect 96777 104147 96805 104175
rect 96839 104147 96867 104175
rect 96901 104147 96929 104175
rect 96963 104147 96991 104175
rect 96777 104085 96805 104113
rect 96839 104085 96867 104113
rect 96901 104085 96929 104113
rect 96963 104085 96991 104113
rect 96777 104023 96805 104051
rect 96839 104023 96867 104051
rect 96901 104023 96929 104051
rect 96963 104023 96991 104051
rect 96777 103961 96805 103989
rect 96839 103961 96867 103989
rect 96901 103961 96929 103989
rect 96963 103961 96991 103989
rect 96777 95147 96805 95175
rect 96839 95147 96867 95175
rect 96901 95147 96929 95175
rect 96963 95147 96991 95175
rect 96777 95085 96805 95113
rect 96839 95085 96867 95113
rect 96901 95085 96929 95113
rect 96963 95085 96991 95113
rect 96777 95023 96805 95051
rect 96839 95023 96867 95051
rect 96901 95023 96929 95051
rect 96963 95023 96991 95051
rect 96777 94961 96805 94989
rect 96839 94961 96867 94989
rect 96901 94961 96929 94989
rect 96963 94961 96991 94989
rect 96777 86147 96805 86175
rect 96839 86147 96867 86175
rect 96901 86147 96929 86175
rect 96963 86147 96991 86175
rect 96777 86085 96805 86113
rect 96839 86085 96867 86113
rect 96901 86085 96929 86113
rect 96963 86085 96991 86113
rect 96777 86023 96805 86051
rect 96839 86023 96867 86051
rect 96901 86023 96929 86051
rect 96963 86023 96991 86051
rect 96777 85961 96805 85989
rect 96839 85961 96867 85989
rect 96901 85961 96929 85989
rect 96963 85961 96991 85989
rect 109939 274961 109967 274989
rect 110001 274961 110029 274989
rect 125299 275147 125327 275175
rect 125361 275147 125389 275175
rect 125299 275085 125327 275113
rect 125361 275085 125389 275113
rect 125299 275023 125327 275051
rect 125361 275023 125389 275051
rect 125299 274961 125327 274989
rect 125361 274961 125389 274989
rect 140659 275147 140687 275175
rect 140721 275147 140749 275175
rect 140659 275085 140687 275113
rect 140721 275085 140749 275113
rect 140659 275023 140687 275051
rect 140721 275023 140749 275051
rect 140659 274961 140687 274989
rect 140721 274961 140749 274989
rect 156019 275147 156047 275175
rect 156081 275147 156109 275175
rect 156019 275085 156047 275113
rect 156081 275085 156109 275113
rect 156019 275023 156047 275051
rect 156081 275023 156109 275051
rect 156019 274961 156047 274989
rect 156081 274961 156109 274989
rect 171379 275147 171407 275175
rect 171441 275147 171469 275175
rect 171379 275085 171407 275113
rect 171441 275085 171469 275113
rect 171379 275023 171407 275051
rect 171441 275023 171469 275051
rect 171379 274961 171407 274989
rect 171441 274961 171469 274989
rect 186739 275147 186767 275175
rect 186801 275147 186829 275175
rect 186739 275085 186767 275113
rect 186801 275085 186829 275113
rect 186739 275023 186767 275051
rect 186801 275023 186829 275051
rect 186739 274961 186767 274989
rect 186801 274961 186829 274989
rect 202099 275147 202127 275175
rect 202161 275147 202189 275175
rect 202099 275085 202127 275113
rect 202161 275085 202189 275113
rect 202099 275023 202127 275051
rect 202161 275023 202189 275051
rect 202099 274961 202127 274989
rect 202161 274961 202189 274989
rect 217459 275147 217487 275175
rect 217521 275147 217549 275175
rect 217459 275085 217487 275113
rect 217521 275085 217549 275113
rect 217459 275023 217487 275051
rect 217521 275023 217549 275051
rect 217459 274961 217487 274989
rect 217521 274961 217549 274989
rect 232819 275147 232847 275175
rect 232881 275147 232909 275175
rect 232819 275085 232847 275113
rect 232881 275085 232909 275113
rect 232819 275023 232847 275051
rect 232881 275023 232909 275051
rect 232819 274961 232847 274989
rect 232881 274961 232909 274989
rect 248179 275147 248207 275175
rect 248241 275147 248269 275175
rect 248179 275085 248207 275113
rect 248241 275085 248269 275113
rect 248179 275023 248207 275051
rect 248241 275023 248269 275051
rect 248179 274961 248207 274989
rect 248241 274961 248269 274989
rect 263539 275147 263567 275175
rect 263601 275147 263629 275175
rect 263539 275085 263567 275113
rect 263601 275085 263629 275113
rect 263539 275023 263567 275051
rect 263601 275023 263629 275051
rect 263539 274961 263567 274989
rect 263601 274961 263629 274989
rect 278899 275147 278927 275175
rect 278961 275147 278989 275175
rect 278899 275085 278927 275113
rect 278961 275085 278989 275113
rect 278899 275023 278927 275051
rect 278961 275023 278989 275051
rect 278899 274961 278927 274989
rect 278961 274961 278989 274989
rect 102259 272147 102287 272175
rect 102321 272147 102349 272175
rect 102259 272085 102287 272113
rect 102321 272085 102349 272113
rect 102259 272023 102287 272051
rect 102321 272023 102349 272051
rect 102259 271961 102287 271989
rect 102321 271961 102349 271989
rect 117619 272147 117647 272175
rect 117681 272147 117709 272175
rect 117619 272085 117647 272113
rect 117681 272085 117709 272113
rect 117619 272023 117647 272051
rect 117681 272023 117709 272051
rect 117619 271961 117647 271989
rect 117681 271961 117709 271989
rect 132979 272147 133007 272175
rect 133041 272147 133069 272175
rect 132979 272085 133007 272113
rect 133041 272085 133069 272113
rect 132979 272023 133007 272051
rect 133041 272023 133069 272051
rect 132979 271961 133007 271989
rect 133041 271961 133069 271989
rect 148339 272147 148367 272175
rect 148401 272147 148429 272175
rect 148339 272085 148367 272113
rect 148401 272085 148429 272113
rect 148339 272023 148367 272051
rect 148401 272023 148429 272051
rect 148339 271961 148367 271989
rect 148401 271961 148429 271989
rect 163699 272147 163727 272175
rect 163761 272147 163789 272175
rect 163699 272085 163727 272113
rect 163761 272085 163789 272113
rect 163699 272023 163727 272051
rect 163761 272023 163789 272051
rect 163699 271961 163727 271989
rect 163761 271961 163789 271989
rect 179059 272147 179087 272175
rect 179121 272147 179149 272175
rect 179059 272085 179087 272113
rect 179121 272085 179149 272113
rect 179059 272023 179087 272051
rect 179121 272023 179149 272051
rect 179059 271961 179087 271989
rect 179121 271961 179149 271989
rect 194419 272147 194447 272175
rect 194481 272147 194509 272175
rect 194419 272085 194447 272113
rect 194481 272085 194509 272113
rect 194419 272023 194447 272051
rect 194481 272023 194509 272051
rect 194419 271961 194447 271989
rect 194481 271961 194509 271989
rect 209779 272147 209807 272175
rect 209841 272147 209869 272175
rect 209779 272085 209807 272113
rect 209841 272085 209869 272113
rect 209779 272023 209807 272051
rect 209841 272023 209869 272051
rect 209779 271961 209807 271989
rect 209841 271961 209869 271989
rect 225139 272147 225167 272175
rect 225201 272147 225229 272175
rect 225139 272085 225167 272113
rect 225201 272085 225229 272113
rect 225139 272023 225167 272051
rect 225201 272023 225229 272051
rect 225139 271961 225167 271989
rect 225201 271961 225229 271989
rect 240499 272147 240527 272175
rect 240561 272147 240589 272175
rect 240499 272085 240527 272113
rect 240561 272085 240589 272113
rect 240499 272023 240527 272051
rect 240561 272023 240589 272051
rect 240499 271961 240527 271989
rect 240561 271961 240589 271989
rect 255859 272147 255887 272175
rect 255921 272147 255949 272175
rect 255859 272085 255887 272113
rect 255921 272085 255949 272113
rect 255859 272023 255887 272051
rect 255921 272023 255949 272051
rect 255859 271961 255887 271989
rect 255921 271961 255949 271989
rect 271219 272147 271247 272175
rect 271281 272147 271309 272175
rect 271219 272085 271247 272113
rect 271281 272085 271309 272113
rect 271219 272023 271247 272051
rect 271281 272023 271309 272051
rect 271219 271961 271247 271989
rect 271281 271961 271309 271989
rect 279237 272147 279265 272175
rect 279299 272147 279327 272175
rect 279361 272147 279389 272175
rect 279423 272147 279451 272175
rect 279237 272085 279265 272113
rect 279299 272085 279327 272113
rect 279361 272085 279389 272113
rect 279423 272085 279451 272113
rect 279237 272023 279265 272051
rect 279299 272023 279327 272051
rect 279361 272023 279389 272051
rect 279423 272023 279451 272051
rect 279237 271961 279265 271989
rect 279299 271961 279327 271989
rect 279361 271961 279389 271989
rect 279423 271961 279451 271989
rect 109939 266147 109967 266175
rect 110001 266147 110029 266175
rect 109939 266085 109967 266113
rect 110001 266085 110029 266113
rect 109939 266023 109967 266051
rect 110001 266023 110029 266051
rect 109939 265961 109967 265989
rect 110001 265961 110029 265989
rect 125299 266147 125327 266175
rect 125361 266147 125389 266175
rect 125299 266085 125327 266113
rect 125361 266085 125389 266113
rect 125299 266023 125327 266051
rect 125361 266023 125389 266051
rect 125299 265961 125327 265989
rect 125361 265961 125389 265989
rect 140659 266147 140687 266175
rect 140721 266147 140749 266175
rect 140659 266085 140687 266113
rect 140721 266085 140749 266113
rect 140659 266023 140687 266051
rect 140721 266023 140749 266051
rect 140659 265961 140687 265989
rect 140721 265961 140749 265989
rect 156019 266147 156047 266175
rect 156081 266147 156109 266175
rect 156019 266085 156047 266113
rect 156081 266085 156109 266113
rect 156019 266023 156047 266051
rect 156081 266023 156109 266051
rect 156019 265961 156047 265989
rect 156081 265961 156109 265989
rect 171379 266147 171407 266175
rect 171441 266147 171469 266175
rect 171379 266085 171407 266113
rect 171441 266085 171469 266113
rect 171379 266023 171407 266051
rect 171441 266023 171469 266051
rect 171379 265961 171407 265989
rect 171441 265961 171469 265989
rect 186739 266147 186767 266175
rect 186801 266147 186829 266175
rect 186739 266085 186767 266113
rect 186801 266085 186829 266113
rect 186739 266023 186767 266051
rect 186801 266023 186829 266051
rect 186739 265961 186767 265989
rect 186801 265961 186829 265989
rect 202099 266147 202127 266175
rect 202161 266147 202189 266175
rect 202099 266085 202127 266113
rect 202161 266085 202189 266113
rect 202099 266023 202127 266051
rect 202161 266023 202189 266051
rect 202099 265961 202127 265989
rect 202161 265961 202189 265989
rect 217459 266147 217487 266175
rect 217521 266147 217549 266175
rect 217459 266085 217487 266113
rect 217521 266085 217549 266113
rect 217459 266023 217487 266051
rect 217521 266023 217549 266051
rect 217459 265961 217487 265989
rect 217521 265961 217549 265989
rect 232819 266147 232847 266175
rect 232881 266147 232909 266175
rect 232819 266085 232847 266113
rect 232881 266085 232909 266113
rect 232819 266023 232847 266051
rect 232881 266023 232909 266051
rect 232819 265961 232847 265989
rect 232881 265961 232909 265989
rect 248179 266147 248207 266175
rect 248241 266147 248269 266175
rect 248179 266085 248207 266113
rect 248241 266085 248269 266113
rect 248179 266023 248207 266051
rect 248241 266023 248269 266051
rect 248179 265961 248207 265989
rect 248241 265961 248269 265989
rect 263539 266147 263567 266175
rect 263601 266147 263629 266175
rect 263539 266085 263567 266113
rect 263601 266085 263629 266113
rect 263539 266023 263567 266051
rect 263601 266023 263629 266051
rect 263539 265961 263567 265989
rect 263601 265961 263629 265989
rect 278899 266147 278927 266175
rect 278961 266147 278989 266175
rect 278899 266085 278927 266113
rect 278961 266085 278989 266113
rect 278899 266023 278927 266051
rect 278961 266023 278989 266051
rect 278899 265961 278927 265989
rect 278961 265961 278989 265989
rect 102259 263147 102287 263175
rect 102321 263147 102349 263175
rect 102259 263085 102287 263113
rect 102321 263085 102349 263113
rect 102259 263023 102287 263051
rect 102321 263023 102349 263051
rect 102259 262961 102287 262989
rect 102321 262961 102349 262989
rect 117619 263147 117647 263175
rect 117681 263147 117709 263175
rect 117619 263085 117647 263113
rect 117681 263085 117709 263113
rect 117619 263023 117647 263051
rect 117681 263023 117709 263051
rect 117619 262961 117647 262989
rect 117681 262961 117709 262989
rect 132979 263147 133007 263175
rect 133041 263147 133069 263175
rect 132979 263085 133007 263113
rect 133041 263085 133069 263113
rect 132979 263023 133007 263051
rect 133041 263023 133069 263051
rect 132979 262961 133007 262989
rect 133041 262961 133069 262989
rect 148339 263147 148367 263175
rect 148401 263147 148429 263175
rect 148339 263085 148367 263113
rect 148401 263085 148429 263113
rect 148339 263023 148367 263051
rect 148401 263023 148429 263051
rect 148339 262961 148367 262989
rect 148401 262961 148429 262989
rect 163699 263147 163727 263175
rect 163761 263147 163789 263175
rect 163699 263085 163727 263113
rect 163761 263085 163789 263113
rect 163699 263023 163727 263051
rect 163761 263023 163789 263051
rect 163699 262961 163727 262989
rect 163761 262961 163789 262989
rect 179059 263147 179087 263175
rect 179121 263147 179149 263175
rect 179059 263085 179087 263113
rect 179121 263085 179149 263113
rect 179059 263023 179087 263051
rect 179121 263023 179149 263051
rect 179059 262961 179087 262989
rect 179121 262961 179149 262989
rect 194419 263147 194447 263175
rect 194481 263147 194509 263175
rect 194419 263085 194447 263113
rect 194481 263085 194509 263113
rect 194419 263023 194447 263051
rect 194481 263023 194509 263051
rect 194419 262961 194447 262989
rect 194481 262961 194509 262989
rect 209779 263147 209807 263175
rect 209841 263147 209869 263175
rect 209779 263085 209807 263113
rect 209841 263085 209869 263113
rect 209779 263023 209807 263051
rect 209841 263023 209869 263051
rect 209779 262961 209807 262989
rect 209841 262961 209869 262989
rect 225139 263147 225167 263175
rect 225201 263147 225229 263175
rect 225139 263085 225167 263113
rect 225201 263085 225229 263113
rect 225139 263023 225167 263051
rect 225201 263023 225229 263051
rect 225139 262961 225167 262989
rect 225201 262961 225229 262989
rect 240499 263147 240527 263175
rect 240561 263147 240589 263175
rect 240499 263085 240527 263113
rect 240561 263085 240589 263113
rect 240499 263023 240527 263051
rect 240561 263023 240589 263051
rect 240499 262961 240527 262989
rect 240561 262961 240589 262989
rect 255859 263147 255887 263175
rect 255921 263147 255949 263175
rect 255859 263085 255887 263113
rect 255921 263085 255949 263113
rect 255859 263023 255887 263051
rect 255921 263023 255949 263051
rect 255859 262961 255887 262989
rect 255921 262961 255949 262989
rect 271219 263147 271247 263175
rect 271281 263147 271309 263175
rect 271219 263085 271247 263113
rect 271281 263085 271309 263113
rect 271219 263023 271247 263051
rect 271281 263023 271309 263051
rect 271219 262961 271247 262989
rect 271281 262961 271309 262989
rect 279237 263147 279265 263175
rect 279299 263147 279327 263175
rect 279361 263147 279389 263175
rect 279423 263147 279451 263175
rect 279237 263085 279265 263113
rect 279299 263085 279327 263113
rect 279361 263085 279389 263113
rect 279423 263085 279451 263113
rect 279237 263023 279265 263051
rect 279299 263023 279327 263051
rect 279361 263023 279389 263051
rect 279423 263023 279451 263051
rect 279237 262961 279265 262989
rect 279299 262961 279327 262989
rect 279361 262961 279389 262989
rect 279423 262961 279451 262989
rect 96777 77147 96805 77175
rect 96839 77147 96867 77175
rect 96901 77147 96929 77175
rect 96963 77147 96991 77175
rect 96777 77085 96805 77113
rect 96839 77085 96867 77113
rect 96901 77085 96929 77113
rect 96963 77085 96991 77113
rect 96777 77023 96805 77051
rect 96839 77023 96867 77051
rect 96901 77023 96929 77051
rect 96963 77023 96991 77051
rect 96777 76961 96805 76989
rect 96839 76961 96867 76989
rect 96901 76961 96929 76989
rect 96963 76961 96991 76989
rect 96777 68147 96805 68175
rect 96839 68147 96867 68175
rect 96901 68147 96929 68175
rect 96963 68147 96991 68175
rect 96777 68085 96805 68113
rect 96839 68085 96867 68113
rect 96901 68085 96929 68113
rect 96963 68085 96991 68113
rect 96777 68023 96805 68051
rect 96839 68023 96867 68051
rect 96901 68023 96929 68051
rect 96963 68023 96991 68051
rect 96777 67961 96805 67989
rect 96839 67961 96867 67989
rect 96901 67961 96929 67989
rect 96963 67961 96991 67989
rect 109939 257147 109967 257175
rect 110001 257147 110029 257175
rect 109939 257085 109967 257113
rect 110001 257085 110029 257113
rect 109939 257023 109967 257051
rect 110001 257023 110029 257051
rect 109939 256961 109967 256989
rect 110001 256961 110029 256989
rect 125299 257147 125327 257175
rect 125361 257147 125389 257175
rect 125299 257085 125327 257113
rect 125361 257085 125389 257113
rect 125299 257023 125327 257051
rect 125361 257023 125389 257051
rect 125299 256961 125327 256989
rect 125361 256961 125389 256989
rect 140659 257147 140687 257175
rect 140721 257147 140749 257175
rect 140659 257085 140687 257113
rect 140721 257085 140749 257113
rect 140659 257023 140687 257051
rect 140721 257023 140749 257051
rect 140659 256961 140687 256989
rect 140721 256961 140749 256989
rect 156019 257147 156047 257175
rect 156081 257147 156109 257175
rect 156019 257085 156047 257113
rect 156081 257085 156109 257113
rect 156019 257023 156047 257051
rect 156081 257023 156109 257051
rect 156019 256961 156047 256989
rect 156081 256961 156109 256989
rect 171379 257147 171407 257175
rect 171441 257147 171469 257175
rect 171379 257085 171407 257113
rect 171441 257085 171469 257113
rect 171379 257023 171407 257051
rect 171441 257023 171469 257051
rect 171379 256961 171407 256989
rect 171441 256961 171469 256989
rect 186739 257147 186767 257175
rect 186801 257147 186829 257175
rect 186739 257085 186767 257113
rect 186801 257085 186829 257113
rect 186739 257023 186767 257051
rect 186801 257023 186829 257051
rect 186739 256961 186767 256989
rect 186801 256961 186829 256989
rect 202099 257147 202127 257175
rect 202161 257147 202189 257175
rect 202099 257085 202127 257113
rect 202161 257085 202189 257113
rect 202099 257023 202127 257051
rect 202161 257023 202189 257051
rect 202099 256961 202127 256989
rect 202161 256961 202189 256989
rect 217459 257147 217487 257175
rect 217521 257147 217549 257175
rect 217459 257085 217487 257113
rect 217521 257085 217549 257113
rect 217459 257023 217487 257051
rect 217521 257023 217549 257051
rect 217459 256961 217487 256989
rect 217521 256961 217549 256989
rect 232819 257147 232847 257175
rect 232881 257147 232909 257175
rect 232819 257085 232847 257113
rect 232881 257085 232909 257113
rect 232819 257023 232847 257051
rect 232881 257023 232909 257051
rect 232819 256961 232847 256989
rect 232881 256961 232909 256989
rect 248179 257147 248207 257175
rect 248241 257147 248269 257175
rect 248179 257085 248207 257113
rect 248241 257085 248269 257113
rect 248179 257023 248207 257051
rect 248241 257023 248269 257051
rect 248179 256961 248207 256989
rect 248241 256961 248269 256989
rect 263539 257147 263567 257175
rect 263601 257147 263629 257175
rect 263539 257085 263567 257113
rect 263601 257085 263629 257113
rect 263539 257023 263567 257051
rect 263601 257023 263629 257051
rect 263539 256961 263567 256989
rect 263601 256961 263629 256989
rect 278899 257147 278927 257175
rect 278961 257147 278989 257175
rect 278899 257085 278927 257113
rect 278961 257085 278989 257113
rect 278899 257023 278927 257051
rect 278961 257023 278989 257051
rect 278899 256961 278927 256989
rect 278961 256961 278989 256989
rect 102259 254147 102287 254175
rect 102321 254147 102349 254175
rect 102259 254085 102287 254113
rect 102321 254085 102349 254113
rect 102259 254023 102287 254051
rect 102321 254023 102349 254051
rect 102259 253961 102287 253989
rect 102321 253961 102349 253989
rect 117619 254147 117647 254175
rect 117681 254147 117709 254175
rect 117619 254085 117647 254113
rect 117681 254085 117709 254113
rect 117619 254023 117647 254051
rect 117681 254023 117709 254051
rect 117619 253961 117647 253989
rect 117681 253961 117709 253989
rect 132979 254147 133007 254175
rect 133041 254147 133069 254175
rect 132979 254085 133007 254113
rect 133041 254085 133069 254113
rect 132979 254023 133007 254051
rect 133041 254023 133069 254051
rect 132979 253961 133007 253989
rect 133041 253961 133069 253989
rect 148339 254147 148367 254175
rect 148401 254147 148429 254175
rect 148339 254085 148367 254113
rect 148401 254085 148429 254113
rect 148339 254023 148367 254051
rect 148401 254023 148429 254051
rect 148339 253961 148367 253989
rect 148401 253961 148429 253989
rect 163699 254147 163727 254175
rect 163761 254147 163789 254175
rect 163699 254085 163727 254113
rect 163761 254085 163789 254113
rect 163699 254023 163727 254051
rect 163761 254023 163789 254051
rect 163699 253961 163727 253989
rect 163761 253961 163789 253989
rect 179059 254147 179087 254175
rect 179121 254147 179149 254175
rect 179059 254085 179087 254113
rect 179121 254085 179149 254113
rect 179059 254023 179087 254051
rect 179121 254023 179149 254051
rect 179059 253961 179087 253989
rect 179121 253961 179149 253989
rect 194419 254147 194447 254175
rect 194481 254147 194509 254175
rect 194419 254085 194447 254113
rect 194481 254085 194509 254113
rect 194419 254023 194447 254051
rect 194481 254023 194509 254051
rect 194419 253961 194447 253989
rect 194481 253961 194509 253989
rect 209779 254147 209807 254175
rect 209841 254147 209869 254175
rect 209779 254085 209807 254113
rect 209841 254085 209869 254113
rect 209779 254023 209807 254051
rect 209841 254023 209869 254051
rect 209779 253961 209807 253989
rect 209841 253961 209869 253989
rect 225139 254147 225167 254175
rect 225201 254147 225229 254175
rect 225139 254085 225167 254113
rect 225201 254085 225229 254113
rect 225139 254023 225167 254051
rect 225201 254023 225229 254051
rect 225139 253961 225167 253989
rect 225201 253961 225229 253989
rect 240499 254147 240527 254175
rect 240561 254147 240589 254175
rect 240499 254085 240527 254113
rect 240561 254085 240589 254113
rect 240499 254023 240527 254051
rect 240561 254023 240589 254051
rect 240499 253961 240527 253989
rect 240561 253961 240589 253989
rect 255859 254147 255887 254175
rect 255921 254147 255949 254175
rect 255859 254085 255887 254113
rect 255921 254085 255949 254113
rect 255859 254023 255887 254051
rect 255921 254023 255949 254051
rect 255859 253961 255887 253989
rect 255921 253961 255949 253989
rect 271219 254147 271247 254175
rect 271281 254147 271309 254175
rect 271219 254085 271247 254113
rect 271281 254085 271309 254113
rect 271219 254023 271247 254051
rect 271281 254023 271309 254051
rect 271219 253961 271247 253989
rect 271281 253961 271309 253989
rect 279237 254147 279265 254175
rect 279299 254147 279327 254175
rect 279361 254147 279389 254175
rect 279423 254147 279451 254175
rect 279237 254085 279265 254113
rect 279299 254085 279327 254113
rect 279361 254085 279389 254113
rect 279423 254085 279451 254113
rect 279237 254023 279265 254051
rect 279299 254023 279327 254051
rect 279361 254023 279389 254051
rect 279423 254023 279451 254051
rect 279237 253961 279265 253989
rect 279299 253961 279327 253989
rect 279361 253961 279389 253989
rect 279423 253961 279451 253989
rect 96777 59147 96805 59175
rect 96839 59147 96867 59175
rect 96901 59147 96929 59175
rect 96963 59147 96991 59175
rect 96777 59085 96805 59113
rect 96839 59085 96867 59113
rect 96901 59085 96929 59113
rect 96963 59085 96991 59113
rect 96777 59023 96805 59051
rect 96839 59023 96867 59051
rect 96901 59023 96929 59051
rect 96963 59023 96991 59051
rect 96777 58961 96805 58989
rect 96839 58961 96867 58989
rect 96901 58961 96929 58989
rect 96963 58961 96991 58989
rect 96777 50147 96805 50175
rect 96839 50147 96867 50175
rect 96901 50147 96929 50175
rect 96963 50147 96991 50175
rect 96777 50085 96805 50113
rect 96839 50085 96867 50113
rect 96901 50085 96929 50113
rect 96963 50085 96991 50113
rect 96777 50023 96805 50051
rect 96839 50023 96867 50051
rect 96901 50023 96929 50051
rect 96963 50023 96991 50051
rect 96777 49961 96805 49989
rect 96839 49961 96867 49989
rect 96901 49961 96929 49989
rect 96963 49961 96991 49989
rect 109939 248147 109967 248175
rect 110001 248147 110029 248175
rect 109939 248085 109967 248113
rect 110001 248085 110029 248113
rect 109939 248023 109967 248051
rect 110001 248023 110029 248051
rect 109939 247961 109967 247989
rect 110001 247961 110029 247989
rect 125299 248147 125327 248175
rect 125361 248147 125389 248175
rect 125299 248085 125327 248113
rect 125361 248085 125389 248113
rect 125299 248023 125327 248051
rect 125361 248023 125389 248051
rect 125299 247961 125327 247989
rect 125361 247961 125389 247989
rect 140659 248147 140687 248175
rect 140721 248147 140749 248175
rect 140659 248085 140687 248113
rect 140721 248085 140749 248113
rect 140659 248023 140687 248051
rect 140721 248023 140749 248051
rect 140659 247961 140687 247989
rect 140721 247961 140749 247989
rect 156019 248147 156047 248175
rect 156081 248147 156109 248175
rect 156019 248085 156047 248113
rect 156081 248085 156109 248113
rect 156019 248023 156047 248051
rect 156081 248023 156109 248051
rect 156019 247961 156047 247989
rect 156081 247961 156109 247989
rect 171379 248147 171407 248175
rect 171441 248147 171469 248175
rect 171379 248085 171407 248113
rect 171441 248085 171469 248113
rect 171379 248023 171407 248051
rect 171441 248023 171469 248051
rect 171379 247961 171407 247989
rect 171441 247961 171469 247989
rect 186739 248147 186767 248175
rect 186801 248147 186829 248175
rect 186739 248085 186767 248113
rect 186801 248085 186829 248113
rect 186739 248023 186767 248051
rect 186801 248023 186829 248051
rect 186739 247961 186767 247989
rect 186801 247961 186829 247989
rect 202099 248147 202127 248175
rect 202161 248147 202189 248175
rect 202099 248085 202127 248113
rect 202161 248085 202189 248113
rect 202099 248023 202127 248051
rect 202161 248023 202189 248051
rect 202099 247961 202127 247989
rect 202161 247961 202189 247989
rect 217459 248147 217487 248175
rect 217521 248147 217549 248175
rect 217459 248085 217487 248113
rect 217521 248085 217549 248113
rect 217459 248023 217487 248051
rect 217521 248023 217549 248051
rect 217459 247961 217487 247989
rect 217521 247961 217549 247989
rect 232819 248147 232847 248175
rect 232881 248147 232909 248175
rect 232819 248085 232847 248113
rect 232881 248085 232909 248113
rect 232819 248023 232847 248051
rect 232881 248023 232909 248051
rect 232819 247961 232847 247989
rect 232881 247961 232909 247989
rect 248179 248147 248207 248175
rect 248241 248147 248269 248175
rect 248179 248085 248207 248113
rect 248241 248085 248269 248113
rect 248179 248023 248207 248051
rect 248241 248023 248269 248051
rect 248179 247961 248207 247989
rect 248241 247961 248269 247989
rect 263539 248147 263567 248175
rect 263601 248147 263629 248175
rect 263539 248085 263567 248113
rect 263601 248085 263629 248113
rect 263539 248023 263567 248051
rect 263601 248023 263629 248051
rect 263539 247961 263567 247989
rect 263601 247961 263629 247989
rect 278899 248147 278927 248175
rect 278961 248147 278989 248175
rect 278899 248085 278927 248113
rect 278961 248085 278989 248113
rect 278899 248023 278927 248051
rect 278961 248023 278989 248051
rect 278899 247961 278927 247989
rect 278961 247961 278989 247989
rect 102259 245147 102287 245175
rect 102321 245147 102349 245175
rect 102259 245085 102287 245113
rect 102321 245085 102349 245113
rect 102259 245023 102287 245051
rect 102321 245023 102349 245051
rect 102259 244961 102287 244989
rect 102321 244961 102349 244989
rect 117619 245147 117647 245175
rect 117681 245147 117709 245175
rect 117619 245085 117647 245113
rect 117681 245085 117709 245113
rect 117619 245023 117647 245051
rect 117681 245023 117709 245051
rect 117619 244961 117647 244989
rect 117681 244961 117709 244989
rect 132979 245147 133007 245175
rect 133041 245147 133069 245175
rect 132979 245085 133007 245113
rect 133041 245085 133069 245113
rect 132979 245023 133007 245051
rect 133041 245023 133069 245051
rect 132979 244961 133007 244989
rect 133041 244961 133069 244989
rect 148339 245147 148367 245175
rect 148401 245147 148429 245175
rect 148339 245085 148367 245113
rect 148401 245085 148429 245113
rect 148339 245023 148367 245051
rect 148401 245023 148429 245051
rect 148339 244961 148367 244989
rect 148401 244961 148429 244989
rect 163699 245147 163727 245175
rect 163761 245147 163789 245175
rect 163699 245085 163727 245113
rect 163761 245085 163789 245113
rect 163699 245023 163727 245051
rect 163761 245023 163789 245051
rect 163699 244961 163727 244989
rect 163761 244961 163789 244989
rect 179059 245147 179087 245175
rect 179121 245147 179149 245175
rect 179059 245085 179087 245113
rect 179121 245085 179149 245113
rect 179059 245023 179087 245051
rect 179121 245023 179149 245051
rect 179059 244961 179087 244989
rect 179121 244961 179149 244989
rect 194419 245147 194447 245175
rect 194481 245147 194509 245175
rect 194419 245085 194447 245113
rect 194481 245085 194509 245113
rect 194419 245023 194447 245051
rect 194481 245023 194509 245051
rect 194419 244961 194447 244989
rect 194481 244961 194509 244989
rect 209779 245147 209807 245175
rect 209841 245147 209869 245175
rect 209779 245085 209807 245113
rect 209841 245085 209869 245113
rect 209779 245023 209807 245051
rect 209841 245023 209869 245051
rect 209779 244961 209807 244989
rect 209841 244961 209869 244989
rect 225139 245147 225167 245175
rect 225201 245147 225229 245175
rect 225139 245085 225167 245113
rect 225201 245085 225229 245113
rect 225139 245023 225167 245051
rect 225201 245023 225229 245051
rect 225139 244961 225167 244989
rect 225201 244961 225229 244989
rect 240499 245147 240527 245175
rect 240561 245147 240589 245175
rect 240499 245085 240527 245113
rect 240561 245085 240589 245113
rect 240499 245023 240527 245051
rect 240561 245023 240589 245051
rect 240499 244961 240527 244989
rect 240561 244961 240589 244989
rect 255859 245147 255887 245175
rect 255921 245147 255949 245175
rect 255859 245085 255887 245113
rect 255921 245085 255949 245113
rect 255859 245023 255887 245051
rect 255921 245023 255949 245051
rect 255859 244961 255887 244989
rect 255921 244961 255949 244989
rect 271219 245147 271247 245175
rect 271281 245147 271309 245175
rect 271219 245085 271247 245113
rect 271281 245085 271309 245113
rect 271219 245023 271247 245051
rect 271281 245023 271309 245051
rect 271219 244961 271247 244989
rect 271281 244961 271309 244989
rect 279237 245147 279265 245175
rect 279299 245147 279327 245175
rect 279361 245147 279389 245175
rect 279423 245147 279451 245175
rect 279237 245085 279265 245113
rect 279299 245085 279327 245113
rect 279361 245085 279389 245113
rect 279423 245085 279451 245113
rect 279237 245023 279265 245051
rect 279299 245023 279327 245051
rect 279361 245023 279389 245051
rect 279423 245023 279451 245051
rect 279237 244961 279265 244989
rect 279299 244961 279327 244989
rect 279361 244961 279389 244989
rect 279423 244961 279451 244989
rect 109939 239147 109967 239175
rect 110001 239147 110029 239175
rect 109939 239085 109967 239113
rect 110001 239085 110029 239113
rect 109939 239023 109967 239051
rect 110001 239023 110029 239051
rect 109939 238961 109967 238989
rect 110001 238961 110029 238989
rect 125299 239147 125327 239175
rect 125361 239147 125389 239175
rect 125299 239085 125327 239113
rect 125361 239085 125389 239113
rect 125299 239023 125327 239051
rect 125361 239023 125389 239051
rect 125299 238961 125327 238989
rect 125361 238961 125389 238989
rect 140659 239147 140687 239175
rect 140721 239147 140749 239175
rect 140659 239085 140687 239113
rect 140721 239085 140749 239113
rect 140659 239023 140687 239051
rect 140721 239023 140749 239051
rect 140659 238961 140687 238989
rect 140721 238961 140749 238989
rect 156019 239147 156047 239175
rect 156081 239147 156109 239175
rect 156019 239085 156047 239113
rect 156081 239085 156109 239113
rect 156019 239023 156047 239051
rect 156081 239023 156109 239051
rect 156019 238961 156047 238989
rect 156081 238961 156109 238989
rect 171379 239147 171407 239175
rect 171441 239147 171469 239175
rect 171379 239085 171407 239113
rect 171441 239085 171469 239113
rect 171379 239023 171407 239051
rect 171441 239023 171469 239051
rect 171379 238961 171407 238989
rect 171441 238961 171469 238989
rect 186739 239147 186767 239175
rect 186801 239147 186829 239175
rect 186739 239085 186767 239113
rect 186801 239085 186829 239113
rect 186739 239023 186767 239051
rect 186801 239023 186829 239051
rect 186739 238961 186767 238989
rect 186801 238961 186829 238989
rect 202099 239147 202127 239175
rect 202161 239147 202189 239175
rect 202099 239085 202127 239113
rect 202161 239085 202189 239113
rect 202099 239023 202127 239051
rect 202161 239023 202189 239051
rect 202099 238961 202127 238989
rect 202161 238961 202189 238989
rect 217459 239147 217487 239175
rect 217521 239147 217549 239175
rect 217459 239085 217487 239113
rect 217521 239085 217549 239113
rect 217459 239023 217487 239051
rect 217521 239023 217549 239051
rect 217459 238961 217487 238989
rect 217521 238961 217549 238989
rect 232819 239147 232847 239175
rect 232881 239147 232909 239175
rect 232819 239085 232847 239113
rect 232881 239085 232909 239113
rect 232819 239023 232847 239051
rect 232881 239023 232909 239051
rect 232819 238961 232847 238989
rect 232881 238961 232909 238989
rect 248179 239147 248207 239175
rect 248241 239147 248269 239175
rect 248179 239085 248207 239113
rect 248241 239085 248269 239113
rect 248179 239023 248207 239051
rect 248241 239023 248269 239051
rect 248179 238961 248207 238989
rect 248241 238961 248269 238989
rect 263539 239147 263567 239175
rect 263601 239147 263629 239175
rect 263539 239085 263567 239113
rect 263601 239085 263629 239113
rect 263539 239023 263567 239051
rect 263601 239023 263629 239051
rect 263539 238961 263567 238989
rect 263601 238961 263629 238989
rect 278899 239147 278927 239175
rect 278961 239147 278989 239175
rect 278899 239085 278927 239113
rect 278961 239085 278989 239113
rect 278899 239023 278927 239051
rect 278961 239023 278989 239051
rect 278899 238961 278927 238989
rect 278961 238961 278989 238989
rect 102259 236147 102287 236175
rect 102321 236147 102349 236175
rect 102259 236085 102287 236113
rect 102321 236085 102349 236113
rect 102259 236023 102287 236051
rect 102321 236023 102349 236051
rect 102259 235961 102287 235989
rect 102321 235961 102349 235989
rect 117619 236147 117647 236175
rect 117681 236147 117709 236175
rect 117619 236085 117647 236113
rect 117681 236085 117709 236113
rect 117619 236023 117647 236051
rect 117681 236023 117709 236051
rect 117619 235961 117647 235989
rect 117681 235961 117709 235989
rect 132979 236147 133007 236175
rect 133041 236147 133069 236175
rect 132979 236085 133007 236113
rect 133041 236085 133069 236113
rect 132979 236023 133007 236051
rect 133041 236023 133069 236051
rect 132979 235961 133007 235989
rect 133041 235961 133069 235989
rect 148339 236147 148367 236175
rect 148401 236147 148429 236175
rect 148339 236085 148367 236113
rect 148401 236085 148429 236113
rect 148339 236023 148367 236051
rect 148401 236023 148429 236051
rect 148339 235961 148367 235989
rect 148401 235961 148429 235989
rect 163699 236147 163727 236175
rect 163761 236147 163789 236175
rect 163699 236085 163727 236113
rect 163761 236085 163789 236113
rect 163699 236023 163727 236051
rect 163761 236023 163789 236051
rect 163699 235961 163727 235989
rect 163761 235961 163789 235989
rect 179059 236147 179087 236175
rect 179121 236147 179149 236175
rect 179059 236085 179087 236113
rect 179121 236085 179149 236113
rect 179059 236023 179087 236051
rect 179121 236023 179149 236051
rect 179059 235961 179087 235989
rect 179121 235961 179149 235989
rect 194419 236147 194447 236175
rect 194481 236147 194509 236175
rect 194419 236085 194447 236113
rect 194481 236085 194509 236113
rect 194419 236023 194447 236051
rect 194481 236023 194509 236051
rect 194419 235961 194447 235989
rect 194481 235961 194509 235989
rect 209779 236147 209807 236175
rect 209841 236147 209869 236175
rect 209779 236085 209807 236113
rect 209841 236085 209869 236113
rect 209779 236023 209807 236051
rect 209841 236023 209869 236051
rect 209779 235961 209807 235989
rect 209841 235961 209869 235989
rect 225139 236147 225167 236175
rect 225201 236147 225229 236175
rect 225139 236085 225167 236113
rect 225201 236085 225229 236113
rect 225139 236023 225167 236051
rect 225201 236023 225229 236051
rect 225139 235961 225167 235989
rect 225201 235961 225229 235989
rect 240499 236147 240527 236175
rect 240561 236147 240589 236175
rect 240499 236085 240527 236113
rect 240561 236085 240589 236113
rect 240499 236023 240527 236051
rect 240561 236023 240589 236051
rect 240499 235961 240527 235989
rect 240561 235961 240589 235989
rect 255859 236147 255887 236175
rect 255921 236147 255949 236175
rect 255859 236085 255887 236113
rect 255921 236085 255949 236113
rect 255859 236023 255887 236051
rect 255921 236023 255949 236051
rect 255859 235961 255887 235989
rect 255921 235961 255949 235989
rect 271219 236147 271247 236175
rect 271281 236147 271309 236175
rect 271219 236085 271247 236113
rect 271281 236085 271309 236113
rect 271219 236023 271247 236051
rect 271281 236023 271309 236051
rect 271219 235961 271247 235989
rect 271281 235961 271309 235989
rect 279237 236147 279265 236175
rect 279299 236147 279327 236175
rect 279361 236147 279389 236175
rect 279423 236147 279451 236175
rect 279237 236085 279265 236113
rect 279299 236085 279327 236113
rect 279361 236085 279389 236113
rect 279423 236085 279451 236113
rect 279237 236023 279265 236051
rect 279299 236023 279327 236051
rect 279361 236023 279389 236051
rect 279423 236023 279451 236051
rect 279237 235961 279265 235989
rect 279299 235961 279327 235989
rect 279361 235961 279389 235989
rect 279423 235961 279451 235989
rect 109939 230147 109967 230175
rect 110001 230147 110029 230175
rect 109939 230085 109967 230113
rect 110001 230085 110029 230113
rect 109939 230023 109967 230051
rect 110001 230023 110029 230051
rect 109939 229961 109967 229989
rect 110001 229961 110029 229989
rect 125299 230147 125327 230175
rect 125361 230147 125389 230175
rect 125299 230085 125327 230113
rect 125361 230085 125389 230113
rect 125299 230023 125327 230051
rect 125361 230023 125389 230051
rect 125299 229961 125327 229989
rect 125361 229961 125389 229989
rect 140659 230147 140687 230175
rect 140721 230147 140749 230175
rect 140659 230085 140687 230113
rect 140721 230085 140749 230113
rect 140659 230023 140687 230051
rect 140721 230023 140749 230051
rect 140659 229961 140687 229989
rect 140721 229961 140749 229989
rect 156019 230147 156047 230175
rect 156081 230147 156109 230175
rect 156019 230085 156047 230113
rect 156081 230085 156109 230113
rect 156019 230023 156047 230051
rect 156081 230023 156109 230051
rect 156019 229961 156047 229989
rect 156081 229961 156109 229989
rect 171379 230147 171407 230175
rect 171441 230147 171469 230175
rect 171379 230085 171407 230113
rect 171441 230085 171469 230113
rect 171379 230023 171407 230051
rect 171441 230023 171469 230051
rect 171379 229961 171407 229989
rect 171441 229961 171469 229989
rect 186739 230147 186767 230175
rect 186801 230147 186829 230175
rect 186739 230085 186767 230113
rect 186801 230085 186829 230113
rect 186739 230023 186767 230051
rect 186801 230023 186829 230051
rect 186739 229961 186767 229989
rect 186801 229961 186829 229989
rect 202099 230147 202127 230175
rect 202161 230147 202189 230175
rect 202099 230085 202127 230113
rect 202161 230085 202189 230113
rect 202099 230023 202127 230051
rect 202161 230023 202189 230051
rect 202099 229961 202127 229989
rect 202161 229961 202189 229989
rect 217459 230147 217487 230175
rect 217521 230147 217549 230175
rect 217459 230085 217487 230113
rect 217521 230085 217549 230113
rect 217459 230023 217487 230051
rect 217521 230023 217549 230051
rect 217459 229961 217487 229989
rect 217521 229961 217549 229989
rect 232819 230147 232847 230175
rect 232881 230147 232909 230175
rect 232819 230085 232847 230113
rect 232881 230085 232909 230113
rect 232819 230023 232847 230051
rect 232881 230023 232909 230051
rect 232819 229961 232847 229989
rect 232881 229961 232909 229989
rect 248179 230147 248207 230175
rect 248241 230147 248269 230175
rect 248179 230085 248207 230113
rect 248241 230085 248269 230113
rect 248179 230023 248207 230051
rect 248241 230023 248269 230051
rect 248179 229961 248207 229989
rect 248241 229961 248269 229989
rect 263539 230147 263567 230175
rect 263601 230147 263629 230175
rect 263539 230085 263567 230113
rect 263601 230085 263629 230113
rect 263539 230023 263567 230051
rect 263601 230023 263629 230051
rect 263539 229961 263567 229989
rect 263601 229961 263629 229989
rect 278899 230147 278927 230175
rect 278961 230147 278989 230175
rect 278899 230085 278927 230113
rect 278961 230085 278989 230113
rect 278899 230023 278927 230051
rect 278961 230023 278989 230051
rect 278899 229961 278927 229989
rect 278961 229961 278989 229989
rect 102259 227147 102287 227175
rect 102321 227147 102349 227175
rect 102259 227085 102287 227113
rect 102321 227085 102349 227113
rect 102259 227023 102287 227051
rect 102321 227023 102349 227051
rect 102259 226961 102287 226989
rect 102321 226961 102349 226989
rect 117619 227147 117647 227175
rect 117681 227147 117709 227175
rect 117619 227085 117647 227113
rect 117681 227085 117709 227113
rect 117619 227023 117647 227051
rect 117681 227023 117709 227051
rect 117619 226961 117647 226989
rect 117681 226961 117709 226989
rect 132979 227147 133007 227175
rect 133041 227147 133069 227175
rect 132979 227085 133007 227113
rect 133041 227085 133069 227113
rect 132979 227023 133007 227051
rect 133041 227023 133069 227051
rect 132979 226961 133007 226989
rect 133041 226961 133069 226989
rect 148339 227147 148367 227175
rect 148401 227147 148429 227175
rect 148339 227085 148367 227113
rect 148401 227085 148429 227113
rect 148339 227023 148367 227051
rect 148401 227023 148429 227051
rect 148339 226961 148367 226989
rect 148401 226961 148429 226989
rect 163699 227147 163727 227175
rect 163761 227147 163789 227175
rect 163699 227085 163727 227113
rect 163761 227085 163789 227113
rect 163699 227023 163727 227051
rect 163761 227023 163789 227051
rect 163699 226961 163727 226989
rect 163761 226961 163789 226989
rect 179059 227147 179087 227175
rect 179121 227147 179149 227175
rect 179059 227085 179087 227113
rect 179121 227085 179149 227113
rect 179059 227023 179087 227051
rect 179121 227023 179149 227051
rect 179059 226961 179087 226989
rect 179121 226961 179149 226989
rect 194419 227147 194447 227175
rect 194481 227147 194509 227175
rect 194419 227085 194447 227113
rect 194481 227085 194509 227113
rect 194419 227023 194447 227051
rect 194481 227023 194509 227051
rect 194419 226961 194447 226989
rect 194481 226961 194509 226989
rect 209779 227147 209807 227175
rect 209841 227147 209869 227175
rect 209779 227085 209807 227113
rect 209841 227085 209869 227113
rect 209779 227023 209807 227051
rect 209841 227023 209869 227051
rect 209779 226961 209807 226989
rect 209841 226961 209869 226989
rect 225139 227147 225167 227175
rect 225201 227147 225229 227175
rect 225139 227085 225167 227113
rect 225201 227085 225229 227113
rect 225139 227023 225167 227051
rect 225201 227023 225229 227051
rect 225139 226961 225167 226989
rect 225201 226961 225229 226989
rect 240499 227147 240527 227175
rect 240561 227147 240589 227175
rect 240499 227085 240527 227113
rect 240561 227085 240589 227113
rect 240499 227023 240527 227051
rect 240561 227023 240589 227051
rect 240499 226961 240527 226989
rect 240561 226961 240589 226989
rect 255859 227147 255887 227175
rect 255921 227147 255949 227175
rect 255859 227085 255887 227113
rect 255921 227085 255949 227113
rect 255859 227023 255887 227051
rect 255921 227023 255949 227051
rect 255859 226961 255887 226989
rect 255921 226961 255949 226989
rect 271219 227147 271247 227175
rect 271281 227147 271309 227175
rect 271219 227085 271247 227113
rect 271281 227085 271309 227113
rect 271219 227023 271247 227051
rect 271281 227023 271309 227051
rect 271219 226961 271247 226989
rect 271281 226961 271309 226989
rect 279237 227147 279265 227175
rect 279299 227147 279327 227175
rect 279361 227147 279389 227175
rect 279423 227147 279451 227175
rect 279237 227085 279265 227113
rect 279299 227085 279327 227113
rect 279361 227085 279389 227113
rect 279423 227085 279451 227113
rect 279237 227023 279265 227051
rect 279299 227023 279327 227051
rect 279361 227023 279389 227051
rect 279423 227023 279451 227051
rect 279237 226961 279265 226989
rect 279299 226961 279327 226989
rect 279361 226961 279389 226989
rect 279423 226961 279451 226989
rect 109939 221147 109967 221175
rect 110001 221147 110029 221175
rect 109939 221085 109967 221113
rect 110001 221085 110029 221113
rect 109939 221023 109967 221051
rect 110001 221023 110029 221051
rect 109939 220961 109967 220989
rect 110001 220961 110029 220989
rect 125299 221147 125327 221175
rect 125361 221147 125389 221175
rect 125299 221085 125327 221113
rect 125361 221085 125389 221113
rect 125299 221023 125327 221051
rect 125361 221023 125389 221051
rect 125299 220961 125327 220989
rect 125361 220961 125389 220989
rect 140659 221147 140687 221175
rect 140721 221147 140749 221175
rect 140659 221085 140687 221113
rect 140721 221085 140749 221113
rect 140659 221023 140687 221051
rect 140721 221023 140749 221051
rect 140659 220961 140687 220989
rect 140721 220961 140749 220989
rect 156019 221147 156047 221175
rect 156081 221147 156109 221175
rect 156019 221085 156047 221113
rect 156081 221085 156109 221113
rect 156019 221023 156047 221051
rect 156081 221023 156109 221051
rect 156019 220961 156047 220989
rect 156081 220961 156109 220989
rect 171379 221147 171407 221175
rect 171441 221147 171469 221175
rect 171379 221085 171407 221113
rect 171441 221085 171469 221113
rect 171379 221023 171407 221051
rect 171441 221023 171469 221051
rect 171379 220961 171407 220989
rect 171441 220961 171469 220989
rect 186739 221147 186767 221175
rect 186801 221147 186829 221175
rect 186739 221085 186767 221113
rect 186801 221085 186829 221113
rect 186739 221023 186767 221051
rect 186801 221023 186829 221051
rect 186739 220961 186767 220989
rect 186801 220961 186829 220989
rect 202099 221147 202127 221175
rect 202161 221147 202189 221175
rect 202099 221085 202127 221113
rect 202161 221085 202189 221113
rect 202099 221023 202127 221051
rect 202161 221023 202189 221051
rect 202099 220961 202127 220989
rect 202161 220961 202189 220989
rect 217459 221147 217487 221175
rect 217521 221147 217549 221175
rect 217459 221085 217487 221113
rect 217521 221085 217549 221113
rect 217459 221023 217487 221051
rect 217521 221023 217549 221051
rect 217459 220961 217487 220989
rect 217521 220961 217549 220989
rect 232819 221147 232847 221175
rect 232881 221147 232909 221175
rect 232819 221085 232847 221113
rect 232881 221085 232909 221113
rect 232819 221023 232847 221051
rect 232881 221023 232909 221051
rect 232819 220961 232847 220989
rect 232881 220961 232909 220989
rect 248179 221147 248207 221175
rect 248241 221147 248269 221175
rect 248179 221085 248207 221113
rect 248241 221085 248269 221113
rect 248179 221023 248207 221051
rect 248241 221023 248269 221051
rect 248179 220961 248207 220989
rect 248241 220961 248269 220989
rect 263539 221147 263567 221175
rect 263601 221147 263629 221175
rect 263539 221085 263567 221113
rect 263601 221085 263629 221113
rect 263539 221023 263567 221051
rect 263601 221023 263629 221051
rect 263539 220961 263567 220989
rect 263601 220961 263629 220989
rect 278899 221147 278927 221175
rect 278961 221147 278989 221175
rect 278899 221085 278927 221113
rect 278961 221085 278989 221113
rect 278899 221023 278927 221051
rect 278961 221023 278989 221051
rect 278899 220961 278927 220989
rect 278961 220961 278989 220989
rect 102259 218147 102287 218175
rect 102321 218147 102349 218175
rect 102259 218085 102287 218113
rect 102321 218085 102349 218113
rect 102259 218023 102287 218051
rect 102321 218023 102349 218051
rect 102259 217961 102287 217989
rect 102321 217961 102349 217989
rect 117619 218147 117647 218175
rect 117681 218147 117709 218175
rect 117619 218085 117647 218113
rect 117681 218085 117709 218113
rect 117619 218023 117647 218051
rect 117681 218023 117709 218051
rect 117619 217961 117647 217989
rect 117681 217961 117709 217989
rect 132979 218147 133007 218175
rect 133041 218147 133069 218175
rect 132979 218085 133007 218113
rect 133041 218085 133069 218113
rect 132979 218023 133007 218051
rect 133041 218023 133069 218051
rect 132979 217961 133007 217989
rect 133041 217961 133069 217989
rect 148339 218147 148367 218175
rect 148401 218147 148429 218175
rect 148339 218085 148367 218113
rect 148401 218085 148429 218113
rect 148339 218023 148367 218051
rect 148401 218023 148429 218051
rect 148339 217961 148367 217989
rect 148401 217961 148429 217989
rect 163699 218147 163727 218175
rect 163761 218147 163789 218175
rect 163699 218085 163727 218113
rect 163761 218085 163789 218113
rect 163699 218023 163727 218051
rect 163761 218023 163789 218051
rect 163699 217961 163727 217989
rect 163761 217961 163789 217989
rect 179059 218147 179087 218175
rect 179121 218147 179149 218175
rect 179059 218085 179087 218113
rect 179121 218085 179149 218113
rect 179059 218023 179087 218051
rect 179121 218023 179149 218051
rect 179059 217961 179087 217989
rect 179121 217961 179149 217989
rect 194419 218147 194447 218175
rect 194481 218147 194509 218175
rect 194419 218085 194447 218113
rect 194481 218085 194509 218113
rect 194419 218023 194447 218051
rect 194481 218023 194509 218051
rect 194419 217961 194447 217989
rect 194481 217961 194509 217989
rect 209779 218147 209807 218175
rect 209841 218147 209869 218175
rect 209779 218085 209807 218113
rect 209841 218085 209869 218113
rect 209779 218023 209807 218051
rect 209841 218023 209869 218051
rect 209779 217961 209807 217989
rect 209841 217961 209869 217989
rect 225139 218147 225167 218175
rect 225201 218147 225229 218175
rect 225139 218085 225167 218113
rect 225201 218085 225229 218113
rect 225139 218023 225167 218051
rect 225201 218023 225229 218051
rect 225139 217961 225167 217989
rect 225201 217961 225229 217989
rect 240499 218147 240527 218175
rect 240561 218147 240589 218175
rect 240499 218085 240527 218113
rect 240561 218085 240589 218113
rect 240499 218023 240527 218051
rect 240561 218023 240589 218051
rect 240499 217961 240527 217989
rect 240561 217961 240589 217989
rect 255859 218147 255887 218175
rect 255921 218147 255949 218175
rect 255859 218085 255887 218113
rect 255921 218085 255949 218113
rect 255859 218023 255887 218051
rect 255921 218023 255949 218051
rect 255859 217961 255887 217989
rect 255921 217961 255949 217989
rect 271219 218147 271247 218175
rect 271281 218147 271309 218175
rect 271219 218085 271247 218113
rect 271281 218085 271309 218113
rect 271219 218023 271247 218051
rect 271281 218023 271309 218051
rect 271219 217961 271247 217989
rect 271281 217961 271309 217989
rect 279237 218147 279265 218175
rect 279299 218147 279327 218175
rect 279361 218147 279389 218175
rect 279423 218147 279451 218175
rect 279237 218085 279265 218113
rect 279299 218085 279327 218113
rect 279361 218085 279389 218113
rect 279423 218085 279451 218113
rect 279237 218023 279265 218051
rect 279299 218023 279327 218051
rect 279361 218023 279389 218051
rect 279423 218023 279451 218051
rect 279237 217961 279265 217989
rect 279299 217961 279327 217989
rect 279361 217961 279389 217989
rect 279423 217961 279451 217989
rect 96777 41147 96805 41175
rect 96839 41147 96867 41175
rect 96901 41147 96929 41175
rect 96963 41147 96991 41175
rect 96777 41085 96805 41113
rect 96839 41085 96867 41113
rect 96901 41085 96929 41113
rect 96963 41085 96991 41113
rect 96777 41023 96805 41051
rect 96839 41023 96867 41051
rect 96901 41023 96929 41051
rect 96963 41023 96991 41051
rect 96777 40961 96805 40989
rect 96839 40961 96867 40989
rect 96901 40961 96929 40989
rect 96963 40961 96991 40989
rect 96777 32147 96805 32175
rect 96839 32147 96867 32175
rect 96901 32147 96929 32175
rect 96963 32147 96991 32175
rect 96777 32085 96805 32113
rect 96839 32085 96867 32113
rect 96901 32085 96929 32113
rect 96963 32085 96991 32113
rect 96777 32023 96805 32051
rect 96839 32023 96867 32051
rect 96901 32023 96929 32051
rect 96963 32023 96991 32051
rect 96777 31961 96805 31989
rect 96839 31961 96867 31989
rect 96901 31961 96929 31989
rect 96963 31961 96991 31989
rect 96777 23147 96805 23175
rect 96839 23147 96867 23175
rect 96901 23147 96929 23175
rect 96963 23147 96991 23175
rect 96777 23085 96805 23113
rect 96839 23085 96867 23113
rect 96901 23085 96929 23113
rect 96963 23085 96991 23113
rect 96777 23023 96805 23051
rect 96839 23023 96867 23051
rect 96901 23023 96929 23051
rect 96963 23023 96991 23051
rect 96777 22961 96805 22989
rect 96839 22961 96867 22989
rect 96901 22961 96929 22989
rect 96963 22961 96991 22989
rect 109939 212147 109967 212175
rect 110001 212147 110029 212175
rect 109939 212085 109967 212113
rect 110001 212085 110029 212113
rect 109939 212023 109967 212051
rect 110001 212023 110029 212051
rect 109939 211961 109967 211989
rect 110001 211961 110029 211989
rect 125299 212147 125327 212175
rect 125361 212147 125389 212175
rect 125299 212085 125327 212113
rect 125361 212085 125389 212113
rect 125299 212023 125327 212051
rect 125361 212023 125389 212051
rect 125299 211961 125327 211989
rect 125361 211961 125389 211989
rect 140659 212147 140687 212175
rect 140721 212147 140749 212175
rect 140659 212085 140687 212113
rect 140721 212085 140749 212113
rect 140659 212023 140687 212051
rect 140721 212023 140749 212051
rect 140659 211961 140687 211989
rect 140721 211961 140749 211989
rect 156019 212147 156047 212175
rect 156081 212147 156109 212175
rect 156019 212085 156047 212113
rect 156081 212085 156109 212113
rect 156019 212023 156047 212051
rect 156081 212023 156109 212051
rect 156019 211961 156047 211989
rect 156081 211961 156109 211989
rect 171379 212147 171407 212175
rect 171441 212147 171469 212175
rect 171379 212085 171407 212113
rect 171441 212085 171469 212113
rect 171379 212023 171407 212051
rect 171441 212023 171469 212051
rect 171379 211961 171407 211989
rect 171441 211961 171469 211989
rect 186739 212147 186767 212175
rect 186801 212147 186829 212175
rect 186739 212085 186767 212113
rect 186801 212085 186829 212113
rect 186739 212023 186767 212051
rect 186801 212023 186829 212051
rect 186739 211961 186767 211989
rect 186801 211961 186829 211989
rect 202099 212147 202127 212175
rect 202161 212147 202189 212175
rect 202099 212085 202127 212113
rect 202161 212085 202189 212113
rect 202099 212023 202127 212051
rect 202161 212023 202189 212051
rect 202099 211961 202127 211989
rect 202161 211961 202189 211989
rect 217459 212147 217487 212175
rect 217521 212147 217549 212175
rect 217459 212085 217487 212113
rect 217521 212085 217549 212113
rect 217459 212023 217487 212051
rect 217521 212023 217549 212051
rect 217459 211961 217487 211989
rect 217521 211961 217549 211989
rect 232819 212147 232847 212175
rect 232881 212147 232909 212175
rect 232819 212085 232847 212113
rect 232881 212085 232909 212113
rect 232819 212023 232847 212051
rect 232881 212023 232909 212051
rect 232819 211961 232847 211989
rect 232881 211961 232909 211989
rect 248179 212147 248207 212175
rect 248241 212147 248269 212175
rect 248179 212085 248207 212113
rect 248241 212085 248269 212113
rect 248179 212023 248207 212051
rect 248241 212023 248269 212051
rect 248179 211961 248207 211989
rect 248241 211961 248269 211989
rect 263539 212147 263567 212175
rect 263601 212147 263629 212175
rect 263539 212085 263567 212113
rect 263601 212085 263629 212113
rect 263539 212023 263567 212051
rect 263601 212023 263629 212051
rect 263539 211961 263567 211989
rect 263601 211961 263629 211989
rect 278899 212147 278927 212175
rect 278961 212147 278989 212175
rect 278899 212085 278927 212113
rect 278961 212085 278989 212113
rect 278899 212023 278927 212051
rect 278961 212023 278989 212051
rect 278899 211961 278927 211989
rect 278961 211961 278989 211989
rect 102259 209147 102287 209175
rect 102321 209147 102349 209175
rect 102259 209085 102287 209113
rect 102321 209085 102349 209113
rect 102259 209023 102287 209051
rect 102321 209023 102349 209051
rect 102259 208961 102287 208989
rect 102321 208961 102349 208989
rect 117619 209147 117647 209175
rect 117681 209147 117709 209175
rect 117619 209085 117647 209113
rect 117681 209085 117709 209113
rect 117619 209023 117647 209051
rect 117681 209023 117709 209051
rect 117619 208961 117647 208989
rect 117681 208961 117709 208989
rect 132979 209147 133007 209175
rect 133041 209147 133069 209175
rect 132979 209085 133007 209113
rect 133041 209085 133069 209113
rect 132979 209023 133007 209051
rect 133041 209023 133069 209051
rect 132979 208961 133007 208989
rect 133041 208961 133069 208989
rect 148339 209147 148367 209175
rect 148401 209147 148429 209175
rect 148339 209085 148367 209113
rect 148401 209085 148429 209113
rect 148339 209023 148367 209051
rect 148401 209023 148429 209051
rect 148339 208961 148367 208989
rect 148401 208961 148429 208989
rect 163699 209147 163727 209175
rect 163761 209147 163789 209175
rect 163699 209085 163727 209113
rect 163761 209085 163789 209113
rect 163699 209023 163727 209051
rect 163761 209023 163789 209051
rect 163699 208961 163727 208989
rect 163761 208961 163789 208989
rect 179059 209147 179087 209175
rect 179121 209147 179149 209175
rect 179059 209085 179087 209113
rect 179121 209085 179149 209113
rect 179059 209023 179087 209051
rect 179121 209023 179149 209051
rect 179059 208961 179087 208989
rect 179121 208961 179149 208989
rect 194419 209147 194447 209175
rect 194481 209147 194509 209175
rect 194419 209085 194447 209113
rect 194481 209085 194509 209113
rect 194419 209023 194447 209051
rect 194481 209023 194509 209051
rect 194419 208961 194447 208989
rect 194481 208961 194509 208989
rect 209779 209147 209807 209175
rect 209841 209147 209869 209175
rect 209779 209085 209807 209113
rect 209841 209085 209869 209113
rect 209779 209023 209807 209051
rect 209841 209023 209869 209051
rect 209779 208961 209807 208989
rect 209841 208961 209869 208989
rect 225139 209147 225167 209175
rect 225201 209147 225229 209175
rect 225139 209085 225167 209113
rect 225201 209085 225229 209113
rect 225139 209023 225167 209051
rect 225201 209023 225229 209051
rect 225139 208961 225167 208989
rect 225201 208961 225229 208989
rect 240499 209147 240527 209175
rect 240561 209147 240589 209175
rect 240499 209085 240527 209113
rect 240561 209085 240589 209113
rect 240499 209023 240527 209051
rect 240561 209023 240589 209051
rect 240499 208961 240527 208989
rect 240561 208961 240589 208989
rect 255859 209147 255887 209175
rect 255921 209147 255949 209175
rect 255859 209085 255887 209113
rect 255921 209085 255949 209113
rect 255859 209023 255887 209051
rect 255921 209023 255949 209051
rect 255859 208961 255887 208989
rect 255921 208961 255949 208989
rect 271219 209147 271247 209175
rect 271281 209147 271309 209175
rect 271219 209085 271247 209113
rect 271281 209085 271309 209113
rect 271219 209023 271247 209051
rect 271281 209023 271309 209051
rect 271219 208961 271247 208989
rect 271281 208961 271309 208989
rect 279237 209147 279265 209175
rect 279299 209147 279327 209175
rect 279361 209147 279389 209175
rect 279423 209147 279451 209175
rect 279237 209085 279265 209113
rect 279299 209085 279327 209113
rect 279361 209085 279389 209113
rect 279423 209085 279451 209113
rect 279237 209023 279265 209051
rect 279299 209023 279327 209051
rect 279361 209023 279389 209051
rect 279423 209023 279451 209051
rect 279237 208961 279265 208989
rect 279299 208961 279327 208989
rect 279361 208961 279389 208989
rect 279423 208961 279451 208989
rect 109939 203147 109967 203175
rect 110001 203147 110029 203175
rect 109939 203085 109967 203113
rect 110001 203085 110029 203113
rect 109939 203023 109967 203051
rect 110001 203023 110029 203051
rect 109939 202961 109967 202989
rect 110001 202961 110029 202989
rect 125299 203147 125327 203175
rect 125361 203147 125389 203175
rect 125299 203085 125327 203113
rect 125361 203085 125389 203113
rect 125299 203023 125327 203051
rect 125361 203023 125389 203051
rect 125299 202961 125327 202989
rect 125361 202961 125389 202989
rect 140659 203147 140687 203175
rect 140721 203147 140749 203175
rect 140659 203085 140687 203113
rect 140721 203085 140749 203113
rect 140659 203023 140687 203051
rect 140721 203023 140749 203051
rect 140659 202961 140687 202989
rect 140721 202961 140749 202989
rect 156019 203147 156047 203175
rect 156081 203147 156109 203175
rect 156019 203085 156047 203113
rect 156081 203085 156109 203113
rect 156019 203023 156047 203051
rect 156081 203023 156109 203051
rect 156019 202961 156047 202989
rect 156081 202961 156109 202989
rect 171379 203147 171407 203175
rect 171441 203147 171469 203175
rect 171379 203085 171407 203113
rect 171441 203085 171469 203113
rect 171379 203023 171407 203051
rect 171441 203023 171469 203051
rect 171379 202961 171407 202989
rect 171441 202961 171469 202989
rect 186739 203147 186767 203175
rect 186801 203147 186829 203175
rect 186739 203085 186767 203113
rect 186801 203085 186829 203113
rect 186739 203023 186767 203051
rect 186801 203023 186829 203051
rect 186739 202961 186767 202989
rect 186801 202961 186829 202989
rect 202099 203147 202127 203175
rect 202161 203147 202189 203175
rect 202099 203085 202127 203113
rect 202161 203085 202189 203113
rect 202099 203023 202127 203051
rect 202161 203023 202189 203051
rect 202099 202961 202127 202989
rect 202161 202961 202189 202989
rect 217459 203147 217487 203175
rect 217521 203147 217549 203175
rect 217459 203085 217487 203113
rect 217521 203085 217549 203113
rect 217459 203023 217487 203051
rect 217521 203023 217549 203051
rect 217459 202961 217487 202989
rect 217521 202961 217549 202989
rect 232819 203147 232847 203175
rect 232881 203147 232909 203175
rect 232819 203085 232847 203113
rect 232881 203085 232909 203113
rect 232819 203023 232847 203051
rect 232881 203023 232909 203051
rect 232819 202961 232847 202989
rect 232881 202961 232909 202989
rect 248179 203147 248207 203175
rect 248241 203147 248269 203175
rect 248179 203085 248207 203113
rect 248241 203085 248269 203113
rect 248179 203023 248207 203051
rect 248241 203023 248269 203051
rect 248179 202961 248207 202989
rect 248241 202961 248269 202989
rect 263539 203147 263567 203175
rect 263601 203147 263629 203175
rect 263539 203085 263567 203113
rect 263601 203085 263629 203113
rect 263539 203023 263567 203051
rect 263601 203023 263629 203051
rect 263539 202961 263567 202989
rect 263601 202961 263629 202989
rect 278899 203147 278927 203175
rect 278961 203147 278989 203175
rect 278899 203085 278927 203113
rect 278961 203085 278989 203113
rect 278899 203023 278927 203051
rect 278961 203023 278989 203051
rect 278899 202961 278927 202989
rect 278961 202961 278989 202989
rect 102259 200147 102287 200175
rect 102321 200147 102349 200175
rect 102259 200085 102287 200113
rect 102321 200085 102349 200113
rect 102259 200023 102287 200051
rect 102321 200023 102349 200051
rect 102259 199961 102287 199989
rect 102321 199961 102349 199989
rect 117619 200147 117647 200175
rect 117681 200147 117709 200175
rect 117619 200085 117647 200113
rect 117681 200085 117709 200113
rect 117619 200023 117647 200051
rect 117681 200023 117709 200051
rect 117619 199961 117647 199989
rect 117681 199961 117709 199989
rect 132979 200147 133007 200175
rect 133041 200147 133069 200175
rect 132979 200085 133007 200113
rect 133041 200085 133069 200113
rect 132979 200023 133007 200051
rect 133041 200023 133069 200051
rect 132979 199961 133007 199989
rect 133041 199961 133069 199989
rect 148339 200147 148367 200175
rect 148401 200147 148429 200175
rect 148339 200085 148367 200113
rect 148401 200085 148429 200113
rect 148339 200023 148367 200051
rect 148401 200023 148429 200051
rect 148339 199961 148367 199989
rect 148401 199961 148429 199989
rect 163699 200147 163727 200175
rect 163761 200147 163789 200175
rect 163699 200085 163727 200113
rect 163761 200085 163789 200113
rect 163699 200023 163727 200051
rect 163761 200023 163789 200051
rect 163699 199961 163727 199989
rect 163761 199961 163789 199989
rect 179059 200147 179087 200175
rect 179121 200147 179149 200175
rect 179059 200085 179087 200113
rect 179121 200085 179149 200113
rect 179059 200023 179087 200051
rect 179121 200023 179149 200051
rect 179059 199961 179087 199989
rect 179121 199961 179149 199989
rect 194419 200147 194447 200175
rect 194481 200147 194509 200175
rect 194419 200085 194447 200113
rect 194481 200085 194509 200113
rect 194419 200023 194447 200051
rect 194481 200023 194509 200051
rect 194419 199961 194447 199989
rect 194481 199961 194509 199989
rect 209779 200147 209807 200175
rect 209841 200147 209869 200175
rect 209779 200085 209807 200113
rect 209841 200085 209869 200113
rect 209779 200023 209807 200051
rect 209841 200023 209869 200051
rect 209779 199961 209807 199989
rect 209841 199961 209869 199989
rect 225139 200147 225167 200175
rect 225201 200147 225229 200175
rect 225139 200085 225167 200113
rect 225201 200085 225229 200113
rect 225139 200023 225167 200051
rect 225201 200023 225229 200051
rect 225139 199961 225167 199989
rect 225201 199961 225229 199989
rect 240499 200147 240527 200175
rect 240561 200147 240589 200175
rect 240499 200085 240527 200113
rect 240561 200085 240589 200113
rect 240499 200023 240527 200051
rect 240561 200023 240589 200051
rect 240499 199961 240527 199989
rect 240561 199961 240589 199989
rect 255859 200147 255887 200175
rect 255921 200147 255949 200175
rect 255859 200085 255887 200113
rect 255921 200085 255949 200113
rect 255859 200023 255887 200051
rect 255921 200023 255949 200051
rect 255859 199961 255887 199989
rect 255921 199961 255949 199989
rect 271219 200147 271247 200175
rect 271281 200147 271309 200175
rect 271219 200085 271247 200113
rect 271281 200085 271309 200113
rect 271219 200023 271247 200051
rect 271281 200023 271309 200051
rect 271219 199961 271247 199989
rect 271281 199961 271309 199989
rect 279237 200147 279265 200175
rect 279299 200147 279327 200175
rect 279361 200147 279389 200175
rect 279423 200147 279451 200175
rect 279237 200085 279265 200113
rect 279299 200085 279327 200113
rect 279361 200085 279389 200113
rect 279423 200085 279451 200113
rect 279237 200023 279265 200051
rect 279299 200023 279327 200051
rect 279361 200023 279389 200051
rect 279423 200023 279451 200051
rect 279237 199961 279265 199989
rect 279299 199961 279327 199989
rect 279361 199961 279389 199989
rect 279423 199961 279451 199989
rect 109939 194147 109967 194175
rect 110001 194147 110029 194175
rect 109939 194085 109967 194113
rect 110001 194085 110029 194113
rect 109939 194023 109967 194051
rect 110001 194023 110029 194051
rect 109939 193961 109967 193989
rect 110001 193961 110029 193989
rect 125299 194147 125327 194175
rect 125361 194147 125389 194175
rect 125299 194085 125327 194113
rect 125361 194085 125389 194113
rect 125299 194023 125327 194051
rect 125361 194023 125389 194051
rect 125299 193961 125327 193989
rect 125361 193961 125389 193989
rect 140659 194147 140687 194175
rect 140721 194147 140749 194175
rect 140659 194085 140687 194113
rect 140721 194085 140749 194113
rect 140659 194023 140687 194051
rect 140721 194023 140749 194051
rect 140659 193961 140687 193989
rect 140721 193961 140749 193989
rect 156019 194147 156047 194175
rect 156081 194147 156109 194175
rect 156019 194085 156047 194113
rect 156081 194085 156109 194113
rect 156019 194023 156047 194051
rect 156081 194023 156109 194051
rect 156019 193961 156047 193989
rect 156081 193961 156109 193989
rect 171379 194147 171407 194175
rect 171441 194147 171469 194175
rect 171379 194085 171407 194113
rect 171441 194085 171469 194113
rect 171379 194023 171407 194051
rect 171441 194023 171469 194051
rect 171379 193961 171407 193989
rect 171441 193961 171469 193989
rect 186739 194147 186767 194175
rect 186801 194147 186829 194175
rect 186739 194085 186767 194113
rect 186801 194085 186829 194113
rect 186739 194023 186767 194051
rect 186801 194023 186829 194051
rect 186739 193961 186767 193989
rect 186801 193961 186829 193989
rect 202099 194147 202127 194175
rect 202161 194147 202189 194175
rect 202099 194085 202127 194113
rect 202161 194085 202189 194113
rect 202099 194023 202127 194051
rect 202161 194023 202189 194051
rect 202099 193961 202127 193989
rect 202161 193961 202189 193989
rect 217459 194147 217487 194175
rect 217521 194147 217549 194175
rect 217459 194085 217487 194113
rect 217521 194085 217549 194113
rect 217459 194023 217487 194051
rect 217521 194023 217549 194051
rect 217459 193961 217487 193989
rect 217521 193961 217549 193989
rect 232819 194147 232847 194175
rect 232881 194147 232909 194175
rect 232819 194085 232847 194113
rect 232881 194085 232909 194113
rect 232819 194023 232847 194051
rect 232881 194023 232909 194051
rect 232819 193961 232847 193989
rect 232881 193961 232909 193989
rect 248179 194147 248207 194175
rect 248241 194147 248269 194175
rect 248179 194085 248207 194113
rect 248241 194085 248269 194113
rect 248179 194023 248207 194051
rect 248241 194023 248269 194051
rect 248179 193961 248207 193989
rect 248241 193961 248269 193989
rect 263539 194147 263567 194175
rect 263601 194147 263629 194175
rect 263539 194085 263567 194113
rect 263601 194085 263629 194113
rect 263539 194023 263567 194051
rect 263601 194023 263629 194051
rect 263539 193961 263567 193989
rect 263601 193961 263629 193989
rect 278899 194147 278927 194175
rect 278961 194147 278989 194175
rect 278899 194085 278927 194113
rect 278961 194085 278989 194113
rect 278899 194023 278927 194051
rect 278961 194023 278989 194051
rect 278899 193961 278927 193989
rect 278961 193961 278989 193989
rect 102259 191147 102287 191175
rect 102321 191147 102349 191175
rect 102259 191085 102287 191113
rect 102321 191085 102349 191113
rect 102259 191023 102287 191051
rect 102321 191023 102349 191051
rect 102259 190961 102287 190989
rect 102321 190961 102349 190989
rect 117619 191147 117647 191175
rect 117681 191147 117709 191175
rect 117619 191085 117647 191113
rect 117681 191085 117709 191113
rect 117619 191023 117647 191051
rect 117681 191023 117709 191051
rect 117619 190961 117647 190989
rect 117681 190961 117709 190989
rect 132979 191147 133007 191175
rect 133041 191147 133069 191175
rect 132979 191085 133007 191113
rect 133041 191085 133069 191113
rect 132979 191023 133007 191051
rect 133041 191023 133069 191051
rect 132979 190961 133007 190989
rect 133041 190961 133069 190989
rect 148339 191147 148367 191175
rect 148401 191147 148429 191175
rect 148339 191085 148367 191113
rect 148401 191085 148429 191113
rect 148339 191023 148367 191051
rect 148401 191023 148429 191051
rect 148339 190961 148367 190989
rect 148401 190961 148429 190989
rect 163699 191147 163727 191175
rect 163761 191147 163789 191175
rect 163699 191085 163727 191113
rect 163761 191085 163789 191113
rect 163699 191023 163727 191051
rect 163761 191023 163789 191051
rect 163699 190961 163727 190989
rect 163761 190961 163789 190989
rect 179059 191147 179087 191175
rect 179121 191147 179149 191175
rect 179059 191085 179087 191113
rect 179121 191085 179149 191113
rect 179059 191023 179087 191051
rect 179121 191023 179149 191051
rect 179059 190961 179087 190989
rect 179121 190961 179149 190989
rect 194419 191147 194447 191175
rect 194481 191147 194509 191175
rect 194419 191085 194447 191113
rect 194481 191085 194509 191113
rect 194419 191023 194447 191051
rect 194481 191023 194509 191051
rect 194419 190961 194447 190989
rect 194481 190961 194509 190989
rect 209779 191147 209807 191175
rect 209841 191147 209869 191175
rect 209779 191085 209807 191113
rect 209841 191085 209869 191113
rect 209779 191023 209807 191051
rect 209841 191023 209869 191051
rect 209779 190961 209807 190989
rect 209841 190961 209869 190989
rect 225139 191147 225167 191175
rect 225201 191147 225229 191175
rect 225139 191085 225167 191113
rect 225201 191085 225229 191113
rect 225139 191023 225167 191051
rect 225201 191023 225229 191051
rect 225139 190961 225167 190989
rect 225201 190961 225229 190989
rect 240499 191147 240527 191175
rect 240561 191147 240589 191175
rect 240499 191085 240527 191113
rect 240561 191085 240589 191113
rect 240499 191023 240527 191051
rect 240561 191023 240589 191051
rect 240499 190961 240527 190989
rect 240561 190961 240589 190989
rect 255859 191147 255887 191175
rect 255921 191147 255949 191175
rect 255859 191085 255887 191113
rect 255921 191085 255949 191113
rect 255859 191023 255887 191051
rect 255921 191023 255949 191051
rect 255859 190961 255887 190989
rect 255921 190961 255949 190989
rect 271219 191147 271247 191175
rect 271281 191147 271309 191175
rect 271219 191085 271247 191113
rect 271281 191085 271309 191113
rect 271219 191023 271247 191051
rect 271281 191023 271309 191051
rect 271219 190961 271247 190989
rect 271281 190961 271309 190989
rect 279237 191147 279265 191175
rect 279299 191147 279327 191175
rect 279361 191147 279389 191175
rect 279423 191147 279451 191175
rect 279237 191085 279265 191113
rect 279299 191085 279327 191113
rect 279361 191085 279389 191113
rect 279423 191085 279451 191113
rect 279237 191023 279265 191051
rect 279299 191023 279327 191051
rect 279361 191023 279389 191051
rect 279423 191023 279451 191051
rect 279237 190961 279265 190989
rect 279299 190961 279327 190989
rect 279361 190961 279389 190989
rect 279423 190961 279451 190989
rect 109939 185147 109967 185175
rect 110001 185147 110029 185175
rect 109939 185085 109967 185113
rect 110001 185085 110029 185113
rect 109939 185023 109967 185051
rect 110001 185023 110029 185051
rect 109939 184961 109967 184989
rect 110001 184961 110029 184989
rect 125299 185147 125327 185175
rect 125361 185147 125389 185175
rect 125299 185085 125327 185113
rect 125361 185085 125389 185113
rect 125299 185023 125327 185051
rect 125361 185023 125389 185051
rect 125299 184961 125327 184989
rect 125361 184961 125389 184989
rect 140659 185147 140687 185175
rect 140721 185147 140749 185175
rect 140659 185085 140687 185113
rect 140721 185085 140749 185113
rect 140659 185023 140687 185051
rect 140721 185023 140749 185051
rect 140659 184961 140687 184989
rect 140721 184961 140749 184989
rect 156019 185147 156047 185175
rect 156081 185147 156109 185175
rect 156019 185085 156047 185113
rect 156081 185085 156109 185113
rect 156019 185023 156047 185051
rect 156081 185023 156109 185051
rect 156019 184961 156047 184989
rect 156081 184961 156109 184989
rect 171379 185147 171407 185175
rect 171441 185147 171469 185175
rect 171379 185085 171407 185113
rect 171441 185085 171469 185113
rect 171379 185023 171407 185051
rect 171441 185023 171469 185051
rect 171379 184961 171407 184989
rect 171441 184961 171469 184989
rect 186739 185147 186767 185175
rect 186801 185147 186829 185175
rect 186739 185085 186767 185113
rect 186801 185085 186829 185113
rect 186739 185023 186767 185051
rect 186801 185023 186829 185051
rect 186739 184961 186767 184989
rect 186801 184961 186829 184989
rect 202099 185147 202127 185175
rect 202161 185147 202189 185175
rect 202099 185085 202127 185113
rect 202161 185085 202189 185113
rect 202099 185023 202127 185051
rect 202161 185023 202189 185051
rect 202099 184961 202127 184989
rect 202161 184961 202189 184989
rect 217459 185147 217487 185175
rect 217521 185147 217549 185175
rect 217459 185085 217487 185113
rect 217521 185085 217549 185113
rect 217459 185023 217487 185051
rect 217521 185023 217549 185051
rect 217459 184961 217487 184989
rect 217521 184961 217549 184989
rect 232819 185147 232847 185175
rect 232881 185147 232909 185175
rect 232819 185085 232847 185113
rect 232881 185085 232909 185113
rect 232819 185023 232847 185051
rect 232881 185023 232909 185051
rect 232819 184961 232847 184989
rect 232881 184961 232909 184989
rect 248179 185147 248207 185175
rect 248241 185147 248269 185175
rect 248179 185085 248207 185113
rect 248241 185085 248269 185113
rect 248179 185023 248207 185051
rect 248241 185023 248269 185051
rect 248179 184961 248207 184989
rect 248241 184961 248269 184989
rect 263539 185147 263567 185175
rect 263601 185147 263629 185175
rect 263539 185085 263567 185113
rect 263601 185085 263629 185113
rect 263539 185023 263567 185051
rect 263601 185023 263629 185051
rect 263539 184961 263567 184989
rect 263601 184961 263629 184989
rect 278899 185147 278927 185175
rect 278961 185147 278989 185175
rect 278899 185085 278927 185113
rect 278961 185085 278989 185113
rect 278899 185023 278927 185051
rect 278961 185023 278989 185051
rect 278899 184961 278927 184989
rect 278961 184961 278989 184989
rect 102259 182147 102287 182175
rect 102321 182147 102349 182175
rect 102259 182085 102287 182113
rect 102321 182085 102349 182113
rect 102259 182023 102287 182051
rect 102321 182023 102349 182051
rect 102259 181961 102287 181989
rect 102321 181961 102349 181989
rect 117619 182147 117647 182175
rect 117681 182147 117709 182175
rect 117619 182085 117647 182113
rect 117681 182085 117709 182113
rect 117619 182023 117647 182051
rect 117681 182023 117709 182051
rect 117619 181961 117647 181989
rect 117681 181961 117709 181989
rect 132979 182147 133007 182175
rect 133041 182147 133069 182175
rect 132979 182085 133007 182113
rect 133041 182085 133069 182113
rect 132979 182023 133007 182051
rect 133041 182023 133069 182051
rect 132979 181961 133007 181989
rect 133041 181961 133069 181989
rect 148339 182147 148367 182175
rect 148401 182147 148429 182175
rect 148339 182085 148367 182113
rect 148401 182085 148429 182113
rect 148339 182023 148367 182051
rect 148401 182023 148429 182051
rect 148339 181961 148367 181989
rect 148401 181961 148429 181989
rect 163699 182147 163727 182175
rect 163761 182147 163789 182175
rect 163699 182085 163727 182113
rect 163761 182085 163789 182113
rect 163699 182023 163727 182051
rect 163761 182023 163789 182051
rect 163699 181961 163727 181989
rect 163761 181961 163789 181989
rect 179059 182147 179087 182175
rect 179121 182147 179149 182175
rect 179059 182085 179087 182113
rect 179121 182085 179149 182113
rect 179059 182023 179087 182051
rect 179121 182023 179149 182051
rect 179059 181961 179087 181989
rect 179121 181961 179149 181989
rect 194419 182147 194447 182175
rect 194481 182147 194509 182175
rect 194419 182085 194447 182113
rect 194481 182085 194509 182113
rect 194419 182023 194447 182051
rect 194481 182023 194509 182051
rect 194419 181961 194447 181989
rect 194481 181961 194509 181989
rect 209779 182147 209807 182175
rect 209841 182147 209869 182175
rect 209779 182085 209807 182113
rect 209841 182085 209869 182113
rect 209779 182023 209807 182051
rect 209841 182023 209869 182051
rect 209779 181961 209807 181989
rect 209841 181961 209869 181989
rect 225139 182147 225167 182175
rect 225201 182147 225229 182175
rect 225139 182085 225167 182113
rect 225201 182085 225229 182113
rect 225139 182023 225167 182051
rect 225201 182023 225229 182051
rect 225139 181961 225167 181989
rect 225201 181961 225229 181989
rect 240499 182147 240527 182175
rect 240561 182147 240589 182175
rect 240499 182085 240527 182113
rect 240561 182085 240589 182113
rect 240499 182023 240527 182051
rect 240561 182023 240589 182051
rect 240499 181961 240527 181989
rect 240561 181961 240589 181989
rect 255859 182147 255887 182175
rect 255921 182147 255949 182175
rect 255859 182085 255887 182113
rect 255921 182085 255949 182113
rect 255859 182023 255887 182051
rect 255921 182023 255949 182051
rect 255859 181961 255887 181989
rect 255921 181961 255949 181989
rect 271219 182147 271247 182175
rect 271281 182147 271309 182175
rect 271219 182085 271247 182113
rect 271281 182085 271309 182113
rect 271219 182023 271247 182051
rect 271281 182023 271309 182051
rect 271219 181961 271247 181989
rect 271281 181961 271309 181989
rect 279237 182147 279265 182175
rect 279299 182147 279327 182175
rect 279361 182147 279389 182175
rect 279423 182147 279451 182175
rect 279237 182085 279265 182113
rect 279299 182085 279327 182113
rect 279361 182085 279389 182113
rect 279423 182085 279451 182113
rect 279237 182023 279265 182051
rect 279299 182023 279327 182051
rect 279361 182023 279389 182051
rect 279423 182023 279451 182051
rect 279237 181961 279265 181989
rect 279299 181961 279327 181989
rect 279361 181961 279389 181989
rect 279423 181961 279451 181989
rect 109939 176147 109967 176175
rect 110001 176147 110029 176175
rect 109939 176085 109967 176113
rect 110001 176085 110029 176113
rect 109939 176023 109967 176051
rect 110001 176023 110029 176051
rect 109939 175961 109967 175989
rect 110001 175961 110029 175989
rect 125299 176147 125327 176175
rect 125361 176147 125389 176175
rect 125299 176085 125327 176113
rect 125361 176085 125389 176113
rect 125299 176023 125327 176051
rect 125361 176023 125389 176051
rect 125299 175961 125327 175989
rect 125361 175961 125389 175989
rect 140659 176147 140687 176175
rect 140721 176147 140749 176175
rect 140659 176085 140687 176113
rect 140721 176085 140749 176113
rect 140659 176023 140687 176051
rect 140721 176023 140749 176051
rect 140659 175961 140687 175989
rect 140721 175961 140749 175989
rect 156019 176147 156047 176175
rect 156081 176147 156109 176175
rect 156019 176085 156047 176113
rect 156081 176085 156109 176113
rect 156019 176023 156047 176051
rect 156081 176023 156109 176051
rect 156019 175961 156047 175989
rect 156081 175961 156109 175989
rect 171379 176147 171407 176175
rect 171441 176147 171469 176175
rect 171379 176085 171407 176113
rect 171441 176085 171469 176113
rect 171379 176023 171407 176051
rect 171441 176023 171469 176051
rect 171379 175961 171407 175989
rect 171441 175961 171469 175989
rect 186739 176147 186767 176175
rect 186801 176147 186829 176175
rect 186739 176085 186767 176113
rect 186801 176085 186829 176113
rect 186739 176023 186767 176051
rect 186801 176023 186829 176051
rect 186739 175961 186767 175989
rect 186801 175961 186829 175989
rect 202099 176147 202127 176175
rect 202161 176147 202189 176175
rect 202099 176085 202127 176113
rect 202161 176085 202189 176113
rect 202099 176023 202127 176051
rect 202161 176023 202189 176051
rect 202099 175961 202127 175989
rect 202161 175961 202189 175989
rect 217459 176147 217487 176175
rect 217521 176147 217549 176175
rect 217459 176085 217487 176113
rect 217521 176085 217549 176113
rect 217459 176023 217487 176051
rect 217521 176023 217549 176051
rect 217459 175961 217487 175989
rect 217521 175961 217549 175989
rect 232819 176147 232847 176175
rect 232881 176147 232909 176175
rect 232819 176085 232847 176113
rect 232881 176085 232909 176113
rect 232819 176023 232847 176051
rect 232881 176023 232909 176051
rect 232819 175961 232847 175989
rect 232881 175961 232909 175989
rect 248179 176147 248207 176175
rect 248241 176147 248269 176175
rect 248179 176085 248207 176113
rect 248241 176085 248269 176113
rect 248179 176023 248207 176051
rect 248241 176023 248269 176051
rect 248179 175961 248207 175989
rect 248241 175961 248269 175989
rect 263539 176147 263567 176175
rect 263601 176147 263629 176175
rect 263539 176085 263567 176113
rect 263601 176085 263629 176113
rect 263539 176023 263567 176051
rect 263601 176023 263629 176051
rect 263539 175961 263567 175989
rect 263601 175961 263629 175989
rect 278899 176147 278927 176175
rect 278961 176147 278989 176175
rect 278899 176085 278927 176113
rect 278961 176085 278989 176113
rect 278899 176023 278927 176051
rect 278961 176023 278989 176051
rect 278899 175961 278927 175989
rect 278961 175961 278989 175989
rect 102259 173147 102287 173175
rect 102321 173147 102349 173175
rect 102259 173085 102287 173113
rect 102321 173085 102349 173113
rect 102259 173023 102287 173051
rect 102321 173023 102349 173051
rect 102259 172961 102287 172989
rect 102321 172961 102349 172989
rect 117619 173147 117647 173175
rect 117681 173147 117709 173175
rect 117619 173085 117647 173113
rect 117681 173085 117709 173113
rect 117619 173023 117647 173051
rect 117681 173023 117709 173051
rect 117619 172961 117647 172989
rect 117681 172961 117709 172989
rect 132979 173147 133007 173175
rect 133041 173147 133069 173175
rect 132979 173085 133007 173113
rect 133041 173085 133069 173113
rect 132979 173023 133007 173051
rect 133041 173023 133069 173051
rect 132979 172961 133007 172989
rect 133041 172961 133069 172989
rect 148339 173147 148367 173175
rect 148401 173147 148429 173175
rect 148339 173085 148367 173113
rect 148401 173085 148429 173113
rect 148339 173023 148367 173051
rect 148401 173023 148429 173051
rect 148339 172961 148367 172989
rect 148401 172961 148429 172989
rect 163699 173147 163727 173175
rect 163761 173147 163789 173175
rect 163699 173085 163727 173113
rect 163761 173085 163789 173113
rect 163699 173023 163727 173051
rect 163761 173023 163789 173051
rect 163699 172961 163727 172989
rect 163761 172961 163789 172989
rect 179059 173147 179087 173175
rect 179121 173147 179149 173175
rect 179059 173085 179087 173113
rect 179121 173085 179149 173113
rect 179059 173023 179087 173051
rect 179121 173023 179149 173051
rect 179059 172961 179087 172989
rect 179121 172961 179149 172989
rect 194419 173147 194447 173175
rect 194481 173147 194509 173175
rect 194419 173085 194447 173113
rect 194481 173085 194509 173113
rect 194419 173023 194447 173051
rect 194481 173023 194509 173051
rect 194419 172961 194447 172989
rect 194481 172961 194509 172989
rect 209779 173147 209807 173175
rect 209841 173147 209869 173175
rect 209779 173085 209807 173113
rect 209841 173085 209869 173113
rect 209779 173023 209807 173051
rect 209841 173023 209869 173051
rect 209779 172961 209807 172989
rect 209841 172961 209869 172989
rect 225139 173147 225167 173175
rect 225201 173147 225229 173175
rect 225139 173085 225167 173113
rect 225201 173085 225229 173113
rect 225139 173023 225167 173051
rect 225201 173023 225229 173051
rect 225139 172961 225167 172989
rect 225201 172961 225229 172989
rect 240499 173147 240527 173175
rect 240561 173147 240589 173175
rect 240499 173085 240527 173113
rect 240561 173085 240589 173113
rect 240499 173023 240527 173051
rect 240561 173023 240589 173051
rect 240499 172961 240527 172989
rect 240561 172961 240589 172989
rect 255859 173147 255887 173175
rect 255921 173147 255949 173175
rect 255859 173085 255887 173113
rect 255921 173085 255949 173113
rect 255859 173023 255887 173051
rect 255921 173023 255949 173051
rect 255859 172961 255887 172989
rect 255921 172961 255949 172989
rect 271219 173147 271247 173175
rect 271281 173147 271309 173175
rect 271219 173085 271247 173113
rect 271281 173085 271309 173113
rect 271219 173023 271247 173051
rect 271281 173023 271309 173051
rect 271219 172961 271247 172989
rect 271281 172961 271309 172989
rect 279237 173147 279265 173175
rect 279299 173147 279327 173175
rect 279361 173147 279389 173175
rect 279423 173147 279451 173175
rect 279237 173085 279265 173113
rect 279299 173085 279327 173113
rect 279361 173085 279389 173113
rect 279423 173085 279451 173113
rect 279237 173023 279265 173051
rect 279299 173023 279327 173051
rect 279361 173023 279389 173051
rect 279423 173023 279451 173051
rect 279237 172961 279265 172989
rect 279299 172961 279327 172989
rect 279361 172961 279389 172989
rect 279423 172961 279451 172989
rect 109939 167147 109967 167175
rect 110001 167147 110029 167175
rect 109939 167085 109967 167113
rect 110001 167085 110029 167113
rect 109939 167023 109967 167051
rect 110001 167023 110029 167051
rect 109939 166961 109967 166989
rect 110001 166961 110029 166989
rect 125299 167147 125327 167175
rect 125361 167147 125389 167175
rect 125299 167085 125327 167113
rect 125361 167085 125389 167113
rect 125299 167023 125327 167051
rect 125361 167023 125389 167051
rect 125299 166961 125327 166989
rect 125361 166961 125389 166989
rect 140659 167147 140687 167175
rect 140721 167147 140749 167175
rect 140659 167085 140687 167113
rect 140721 167085 140749 167113
rect 140659 167023 140687 167051
rect 140721 167023 140749 167051
rect 140659 166961 140687 166989
rect 140721 166961 140749 166989
rect 156019 167147 156047 167175
rect 156081 167147 156109 167175
rect 156019 167085 156047 167113
rect 156081 167085 156109 167113
rect 156019 167023 156047 167051
rect 156081 167023 156109 167051
rect 156019 166961 156047 166989
rect 156081 166961 156109 166989
rect 171379 167147 171407 167175
rect 171441 167147 171469 167175
rect 171379 167085 171407 167113
rect 171441 167085 171469 167113
rect 171379 167023 171407 167051
rect 171441 167023 171469 167051
rect 171379 166961 171407 166989
rect 171441 166961 171469 166989
rect 186739 167147 186767 167175
rect 186801 167147 186829 167175
rect 186739 167085 186767 167113
rect 186801 167085 186829 167113
rect 186739 167023 186767 167051
rect 186801 167023 186829 167051
rect 186739 166961 186767 166989
rect 186801 166961 186829 166989
rect 202099 167147 202127 167175
rect 202161 167147 202189 167175
rect 202099 167085 202127 167113
rect 202161 167085 202189 167113
rect 202099 167023 202127 167051
rect 202161 167023 202189 167051
rect 202099 166961 202127 166989
rect 202161 166961 202189 166989
rect 217459 167147 217487 167175
rect 217521 167147 217549 167175
rect 217459 167085 217487 167113
rect 217521 167085 217549 167113
rect 217459 167023 217487 167051
rect 217521 167023 217549 167051
rect 217459 166961 217487 166989
rect 217521 166961 217549 166989
rect 232819 167147 232847 167175
rect 232881 167147 232909 167175
rect 232819 167085 232847 167113
rect 232881 167085 232909 167113
rect 232819 167023 232847 167051
rect 232881 167023 232909 167051
rect 232819 166961 232847 166989
rect 232881 166961 232909 166989
rect 248179 167147 248207 167175
rect 248241 167147 248269 167175
rect 248179 167085 248207 167113
rect 248241 167085 248269 167113
rect 248179 167023 248207 167051
rect 248241 167023 248269 167051
rect 248179 166961 248207 166989
rect 248241 166961 248269 166989
rect 263539 167147 263567 167175
rect 263601 167147 263629 167175
rect 263539 167085 263567 167113
rect 263601 167085 263629 167113
rect 263539 167023 263567 167051
rect 263601 167023 263629 167051
rect 263539 166961 263567 166989
rect 263601 166961 263629 166989
rect 278899 167147 278927 167175
rect 278961 167147 278989 167175
rect 278899 167085 278927 167113
rect 278961 167085 278989 167113
rect 278899 167023 278927 167051
rect 278961 167023 278989 167051
rect 278899 166961 278927 166989
rect 278961 166961 278989 166989
rect 102259 164147 102287 164175
rect 102321 164147 102349 164175
rect 102259 164085 102287 164113
rect 102321 164085 102349 164113
rect 102259 164023 102287 164051
rect 102321 164023 102349 164051
rect 102259 163961 102287 163989
rect 102321 163961 102349 163989
rect 117619 164147 117647 164175
rect 117681 164147 117709 164175
rect 117619 164085 117647 164113
rect 117681 164085 117709 164113
rect 117619 164023 117647 164051
rect 117681 164023 117709 164051
rect 117619 163961 117647 163989
rect 117681 163961 117709 163989
rect 132979 164147 133007 164175
rect 133041 164147 133069 164175
rect 132979 164085 133007 164113
rect 133041 164085 133069 164113
rect 132979 164023 133007 164051
rect 133041 164023 133069 164051
rect 132979 163961 133007 163989
rect 133041 163961 133069 163989
rect 148339 164147 148367 164175
rect 148401 164147 148429 164175
rect 148339 164085 148367 164113
rect 148401 164085 148429 164113
rect 148339 164023 148367 164051
rect 148401 164023 148429 164051
rect 148339 163961 148367 163989
rect 148401 163961 148429 163989
rect 163699 164147 163727 164175
rect 163761 164147 163789 164175
rect 163699 164085 163727 164113
rect 163761 164085 163789 164113
rect 163699 164023 163727 164051
rect 163761 164023 163789 164051
rect 163699 163961 163727 163989
rect 163761 163961 163789 163989
rect 179059 164147 179087 164175
rect 179121 164147 179149 164175
rect 179059 164085 179087 164113
rect 179121 164085 179149 164113
rect 179059 164023 179087 164051
rect 179121 164023 179149 164051
rect 179059 163961 179087 163989
rect 179121 163961 179149 163989
rect 194419 164147 194447 164175
rect 194481 164147 194509 164175
rect 194419 164085 194447 164113
rect 194481 164085 194509 164113
rect 194419 164023 194447 164051
rect 194481 164023 194509 164051
rect 194419 163961 194447 163989
rect 194481 163961 194509 163989
rect 209779 164147 209807 164175
rect 209841 164147 209869 164175
rect 209779 164085 209807 164113
rect 209841 164085 209869 164113
rect 209779 164023 209807 164051
rect 209841 164023 209869 164051
rect 209779 163961 209807 163989
rect 209841 163961 209869 163989
rect 225139 164147 225167 164175
rect 225201 164147 225229 164175
rect 225139 164085 225167 164113
rect 225201 164085 225229 164113
rect 225139 164023 225167 164051
rect 225201 164023 225229 164051
rect 225139 163961 225167 163989
rect 225201 163961 225229 163989
rect 240499 164147 240527 164175
rect 240561 164147 240589 164175
rect 240499 164085 240527 164113
rect 240561 164085 240589 164113
rect 240499 164023 240527 164051
rect 240561 164023 240589 164051
rect 240499 163961 240527 163989
rect 240561 163961 240589 163989
rect 255859 164147 255887 164175
rect 255921 164147 255949 164175
rect 255859 164085 255887 164113
rect 255921 164085 255949 164113
rect 255859 164023 255887 164051
rect 255921 164023 255949 164051
rect 255859 163961 255887 163989
rect 255921 163961 255949 163989
rect 271219 164147 271247 164175
rect 271281 164147 271309 164175
rect 271219 164085 271247 164113
rect 271281 164085 271309 164113
rect 271219 164023 271247 164051
rect 271281 164023 271309 164051
rect 271219 163961 271247 163989
rect 271281 163961 271309 163989
rect 279237 164147 279265 164175
rect 279299 164147 279327 164175
rect 279361 164147 279389 164175
rect 279423 164147 279451 164175
rect 279237 164085 279265 164113
rect 279299 164085 279327 164113
rect 279361 164085 279389 164113
rect 279423 164085 279451 164113
rect 279237 164023 279265 164051
rect 279299 164023 279327 164051
rect 279361 164023 279389 164051
rect 279423 164023 279451 164051
rect 279237 163961 279265 163989
rect 279299 163961 279327 163989
rect 279361 163961 279389 163989
rect 279423 163961 279451 163989
rect 109939 158147 109967 158175
rect 110001 158147 110029 158175
rect 109939 158085 109967 158113
rect 110001 158085 110029 158113
rect 109939 158023 109967 158051
rect 110001 158023 110029 158051
rect 109939 157961 109967 157989
rect 110001 157961 110029 157989
rect 125299 158147 125327 158175
rect 125361 158147 125389 158175
rect 125299 158085 125327 158113
rect 125361 158085 125389 158113
rect 125299 158023 125327 158051
rect 125361 158023 125389 158051
rect 125299 157961 125327 157989
rect 125361 157961 125389 157989
rect 140659 158147 140687 158175
rect 140721 158147 140749 158175
rect 140659 158085 140687 158113
rect 140721 158085 140749 158113
rect 140659 158023 140687 158051
rect 140721 158023 140749 158051
rect 140659 157961 140687 157989
rect 140721 157961 140749 157989
rect 156019 158147 156047 158175
rect 156081 158147 156109 158175
rect 156019 158085 156047 158113
rect 156081 158085 156109 158113
rect 156019 158023 156047 158051
rect 156081 158023 156109 158051
rect 156019 157961 156047 157989
rect 156081 157961 156109 157989
rect 171379 158147 171407 158175
rect 171441 158147 171469 158175
rect 171379 158085 171407 158113
rect 171441 158085 171469 158113
rect 171379 158023 171407 158051
rect 171441 158023 171469 158051
rect 171379 157961 171407 157989
rect 171441 157961 171469 157989
rect 186739 158147 186767 158175
rect 186801 158147 186829 158175
rect 186739 158085 186767 158113
rect 186801 158085 186829 158113
rect 186739 158023 186767 158051
rect 186801 158023 186829 158051
rect 186739 157961 186767 157989
rect 186801 157961 186829 157989
rect 202099 158147 202127 158175
rect 202161 158147 202189 158175
rect 202099 158085 202127 158113
rect 202161 158085 202189 158113
rect 202099 158023 202127 158051
rect 202161 158023 202189 158051
rect 202099 157961 202127 157989
rect 202161 157961 202189 157989
rect 217459 158147 217487 158175
rect 217521 158147 217549 158175
rect 217459 158085 217487 158113
rect 217521 158085 217549 158113
rect 217459 158023 217487 158051
rect 217521 158023 217549 158051
rect 217459 157961 217487 157989
rect 217521 157961 217549 157989
rect 232819 158147 232847 158175
rect 232881 158147 232909 158175
rect 232819 158085 232847 158113
rect 232881 158085 232909 158113
rect 232819 158023 232847 158051
rect 232881 158023 232909 158051
rect 232819 157961 232847 157989
rect 232881 157961 232909 157989
rect 248179 158147 248207 158175
rect 248241 158147 248269 158175
rect 248179 158085 248207 158113
rect 248241 158085 248269 158113
rect 248179 158023 248207 158051
rect 248241 158023 248269 158051
rect 248179 157961 248207 157989
rect 248241 157961 248269 157989
rect 263539 158147 263567 158175
rect 263601 158147 263629 158175
rect 263539 158085 263567 158113
rect 263601 158085 263629 158113
rect 263539 158023 263567 158051
rect 263601 158023 263629 158051
rect 263539 157961 263567 157989
rect 263601 157961 263629 157989
rect 278899 158147 278927 158175
rect 278961 158147 278989 158175
rect 278899 158085 278927 158113
rect 278961 158085 278989 158113
rect 278899 158023 278927 158051
rect 278961 158023 278989 158051
rect 278899 157961 278927 157989
rect 278961 157961 278989 157989
rect 102259 155147 102287 155175
rect 102321 155147 102349 155175
rect 102259 155085 102287 155113
rect 102321 155085 102349 155113
rect 102259 155023 102287 155051
rect 102321 155023 102349 155051
rect 102259 154961 102287 154989
rect 102321 154961 102349 154989
rect 117619 155147 117647 155175
rect 117681 155147 117709 155175
rect 117619 155085 117647 155113
rect 117681 155085 117709 155113
rect 117619 155023 117647 155051
rect 117681 155023 117709 155051
rect 117619 154961 117647 154989
rect 117681 154961 117709 154989
rect 132979 155147 133007 155175
rect 133041 155147 133069 155175
rect 132979 155085 133007 155113
rect 133041 155085 133069 155113
rect 132979 155023 133007 155051
rect 133041 155023 133069 155051
rect 132979 154961 133007 154989
rect 133041 154961 133069 154989
rect 148339 155147 148367 155175
rect 148401 155147 148429 155175
rect 148339 155085 148367 155113
rect 148401 155085 148429 155113
rect 148339 155023 148367 155051
rect 148401 155023 148429 155051
rect 148339 154961 148367 154989
rect 148401 154961 148429 154989
rect 163699 155147 163727 155175
rect 163761 155147 163789 155175
rect 163699 155085 163727 155113
rect 163761 155085 163789 155113
rect 163699 155023 163727 155051
rect 163761 155023 163789 155051
rect 163699 154961 163727 154989
rect 163761 154961 163789 154989
rect 179059 155147 179087 155175
rect 179121 155147 179149 155175
rect 179059 155085 179087 155113
rect 179121 155085 179149 155113
rect 179059 155023 179087 155051
rect 179121 155023 179149 155051
rect 179059 154961 179087 154989
rect 179121 154961 179149 154989
rect 194419 155147 194447 155175
rect 194481 155147 194509 155175
rect 194419 155085 194447 155113
rect 194481 155085 194509 155113
rect 194419 155023 194447 155051
rect 194481 155023 194509 155051
rect 194419 154961 194447 154989
rect 194481 154961 194509 154989
rect 209779 155147 209807 155175
rect 209841 155147 209869 155175
rect 209779 155085 209807 155113
rect 209841 155085 209869 155113
rect 209779 155023 209807 155051
rect 209841 155023 209869 155051
rect 209779 154961 209807 154989
rect 209841 154961 209869 154989
rect 225139 155147 225167 155175
rect 225201 155147 225229 155175
rect 225139 155085 225167 155113
rect 225201 155085 225229 155113
rect 225139 155023 225167 155051
rect 225201 155023 225229 155051
rect 225139 154961 225167 154989
rect 225201 154961 225229 154989
rect 240499 155147 240527 155175
rect 240561 155147 240589 155175
rect 240499 155085 240527 155113
rect 240561 155085 240589 155113
rect 240499 155023 240527 155051
rect 240561 155023 240589 155051
rect 240499 154961 240527 154989
rect 240561 154961 240589 154989
rect 255859 155147 255887 155175
rect 255921 155147 255949 155175
rect 255859 155085 255887 155113
rect 255921 155085 255949 155113
rect 255859 155023 255887 155051
rect 255921 155023 255949 155051
rect 255859 154961 255887 154989
rect 255921 154961 255949 154989
rect 271219 155147 271247 155175
rect 271281 155147 271309 155175
rect 271219 155085 271247 155113
rect 271281 155085 271309 155113
rect 271219 155023 271247 155051
rect 271281 155023 271309 155051
rect 271219 154961 271247 154989
rect 271281 154961 271309 154989
rect 279237 155147 279265 155175
rect 279299 155147 279327 155175
rect 279361 155147 279389 155175
rect 279423 155147 279451 155175
rect 279237 155085 279265 155113
rect 279299 155085 279327 155113
rect 279361 155085 279389 155113
rect 279423 155085 279451 155113
rect 279237 155023 279265 155051
rect 279299 155023 279327 155051
rect 279361 155023 279389 155051
rect 279423 155023 279451 155051
rect 279237 154961 279265 154989
rect 279299 154961 279327 154989
rect 279361 154961 279389 154989
rect 279423 154961 279451 154989
rect 109939 149147 109967 149175
rect 110001 149147 110029 149175
rect 109939 149085 109967 149113
rect 110001 149085 110029 149113
rect 109939 149023 109967 149051
rect 110001 149023 110029 149051
rect 109939 148961 109967 148989
rect 110001 148961 110029 148989
rect 125299 149147 125327 149175
rect 125361 149147 125389 149175
rect 125299 149085 125327 149113
rect 125361 149085 125389 149113
rect 125299 149023 125327 149051
rect 125361 149023 125389 149051
rect 125299 148961 125327 148989
rect 125361 148961 125389 148989
rect 140659 149147 140687 149175
rect 140721 149147 140749 149175
rect 140659 149085 140687 149113
rect 140721 149085 140749 149113
rect 140659 149023 140687 149051
rect 140721 149023 140749 149051
rect 140659 148961 140687 148989
rect 140721 148961 140749 148989
rect 156019 149147 156047 149175
rect 156081 149147 156109 149175
rect 156019 149085 156047 149113
rect 156081 149085 156109 149113
rect 156019 149023 156047 149051
rect 156081 149023 156109 149051
rect 156019 148961 156047 148989
rect 156081 148961 156109 148989
rect 171379 149147 171407 149175
rect 171441 149147 171469 149175
rect 171379 149085 171407 149113
rect 171441 149085 171469 149113
rect 171379 149023 171407 149051
rect 171441 149023 171469 149051
rect 171379 148961 171407 148989
rect 171441 148961 171469 148989
rect 186739 149147 186767 149175
rect 186801 149147 186829 149175
rect 186739 149085 186767 149113
rect 186801 149085 186829 149113
rect 186739 149023 186767 149051
rect 186801 149023 186829 149051
rect 186739 148961 186767 148989
rect 186801 148961 186829 148989
rect 202099 149147 202127 149175
rect 202161 149147 202189 149175
rect 202099 149085 202127 149113
rect 202161 149085 202189 149113
rect 202099 149023 202127 149051
rect 202161 149023 202189 149051
rect 202099 148961 202127 148989
rect 202161 148961 202189 148989
rect 217459 149147 217487 149175
rect 217521 149147 217549 149175
rect 217459 149085 217487 149113
rect 217521 149085 217549 149113
rect 217459 149023 217487 149051
rect 217521 149023 217549 149051
rect 217459 148961 217487 148989
rect 217521 148961 217549 148989
rect 232819 149147 232847 149175
rect 232881 149147 232909 149175
rect 232819 149085 232847 149113
rect 232881 149085 232909 149113
rect 232819 149023 232847 149051
rect 232881 149023 232909 149051
rect 232819 148961 232847 148989
rect 232881 148961 232909 148989
rect 248179 149147 248207 149175
rect 248241 149147 248269 149175
rect 248179 149085 248207 149113
rect 248241 149085 248269 149113
rect 248179 149023 248207 149051
rect 248241 149023 248269 149051
rect 248179 148961 248207 148989
rect 248241 148961 248269 148989
rect 263539 149147 263567 149175
rect 263601 149147 263629 149175
rect 263539 149085 263567 149113
rect 263601 149085 263629 149113
rect 263539 149023 263567 149051
rect 263601 149023 263629 149051
rect 263539 148961 263567 148989
rect 263601 148961 263629 148989
rect 278899 149147 278927 149175
rect 278961 149147 278989 149175
rect 278899 149085 278927 149113
rect 278961 149085 278989 149113
rect 278899 149023 278927 149051
rect 278961 149023 278989 149051
rect 278899 148961 278927 148989
rect 278961 148961 278989 148989
rect 102259 146147 102287 146175
rect 102321 146147 102349 146175
rect 102259 146085 102287 146113
rect 102321 146085 102349 146113
rect 102259 146023 102287 146051
rect 102321 146023 102349 146051
rect 102259 145961 102287 145989
rect 102321 145961 102349 145989
rect 117619 146147 117647 146175
rect 117681 146147 117709 146175
rect 117619 146085 117647 146113
rect 117681 146085 117709 146113
rect 117619 146023 117647 146051
rect 117681 146023 117709 146051
rect 117619 145961 117647 145989
rect 117681 145961 117709 145989
rect 132979 146147 133007 146175
rect 133041 146147 133069 146175
rect 132979 146085 133007 146113
rect 133041 146085 133069 146113
rect 132979 146023 133007 146051
rect 133041 146023 133069 146051
rect 132979 145961 133007 145989
rect 133041 145961 133069 145989
rect 148339 146147 148367 146175
rect 148401 146147 148429 146175
rect 148339 146085 148367 146113
rect 148401 146085 148429 146113
rect 148339 146023 148367 146051
rect 148401 146023 148429 146051
rect 148339 145961 148367 145989
rect 148401 145961 148429 145989
rect 163699 146147 163727 146175
rect 163761 146147 163789 146175
rect 163699 146085 163727 146113
rect 163761 146085 163789 146113
rect 163699 146023 163727 146051
rect 163761 146023 163789 146051
rect 163699 145961 163727 145989
rect 163761 145961 163789 145989
rect 179059 146147 179087 146175
rect 179121 146147 179149 146175
rect 179059 146085 179087 146113
rect 179121 146085 179149 146113
rect 179059 146023 179087 146051
rect 179121 146023 179149 146051
rect 179059 145961 179087 145989
rect 179121 145961 179149 145989
rect 194419 146147 194447 146175
rect 194481 146147 194509 146175
rect 194419 146085 194447 146113
rect 194481 146085 194509 146113
rect 194419 146023 194447 146051
rect 194481 146023 194509 146051
rect 194419 145961 194447 145989
rect 194481 145961 194509 145989
rect 209779 146147 209807 146175
rect 209841 146147 209869 146175
rect 209779 146085 209807 146113
rect 209841 146085 209869 146113
rect 209779 146023 209807 146051
rect 209841 146023 209869 146051
rect 209779 145961 209807 145989
rect 209841 145961 209869 145989
rect 225139 146147 225167 146175
rect 225201 146147 225229 146175
rect 225139 146085 225167 146113
rect 225201 146085 225229 146113
rect 225139 146023 225167 146051
rect 225201 146023 225229 146051
rect 225139 145961 225167 145989
rect 225201 145961 225229 145989
rect 240499 146147 240527 146175
rect 240561 146147 240589 146175
rect 240499 146085 240527 146113
rect 240561 146085 240589 146113
rect 240499 146023 240527 146051
rect 240561 146023 240589 146051
rect 240499 145961 240527 145989
rect 240561 145961 240589 145989
rect 255859 146147 255887 146175
rect 255921 146147 255949 146175
rect 255859 146085 255887 146113
rect 255921 146085 255949 146113
rect 255859 146023 255887 146051
rect 255921 146023 255949 146051
rect 255859 145961 255887 145989
rect 255921 145961 255949 145989
rect 271219 146147 271247 146175
rect 271281 146147 271309 146175
rect 271219 146085 271247 146113
rect 271281 146085 271309 146113
rect 271219 146023 271247 146051
rect 271281 146023 271309 146051
rect 271219 145961 271247 145989
rect 271281 145961 271309 145989
rect 279237 146147 279265 146175
rect 279299 146147 279327 146175
rect 279361 146147 279389 146175
rect 279423 146147 279451 146175
rect 279237 146085 279265 146113
rect 279299 146085 279327 146113
rect 279361 146085 279389 146113
rect 279423 146085 279451 146113
rect 279237 146023 279265 146051
rect 279299 146023 279327 146051
rect 279361 146023 279389 146051
rect 279423 146023 279451 146051
rect 279237 145961 279265 145989
rect 279299 145961 279327 145989
rect 279361 145961 279389 145989
rect 279423 145961 279451 145989
rect 109939 140147 109967 140175
rect 110001 140147 110029 140175
rect 109939 140085 109967 140113
rect 110001 140085 110029 140113
rect 109939 140023 109967 140051
rect 110001 140023 110029 140051
rect 109939 139961 109967 139989
rect 110001 139961 110029 139989
rect 125299 140147 125327 140175
rect 125361 140147 125389 140175
rect 125299 140085 125327 140113
rect 125361 140085 125389 140113
rect 125299 140023 125327 140051
rect 125361 140023 125389 140051
rect 125299 139961 125327 139989
rect 125361 139961 125389 139989
rect 140659 140147 140687 140175
rect 140721 140147 140749 140175
rect 140659 140085 140687 140113
rect 140721 140085 140749 140113
rect 140659 140023 140687 140051
rect 140721 140023 140749 140051
rect 140659 139961 140687 139989
rect 140721 139961 140749 139989
rect 156019 140147 156047 140175
rect 156081 140147 156109 140175
rect 156019 140085 156047 140113
rect 156081 140085 156109 140113
rect 156019 140023 156047 140051
rect 156081 140023 156109 140051
rect 156019 139961 156047 139989
rect 156081 139961 156109 139989
rect 171379 140147 171407 140175
rect 171441 140147 171469 140175
rect 171379 140085 171407 140113
rect 171441 140085 171469 140113
rect 171379 140023 171407 140051
rect 171441 140023 171469 140051
rect 171379 139961 171407 139989
rect 171441 139961 171469 139989
rect 186739 140147 186767 140175
rect 186801 140147 186829 140175
rect 186739 140085 186767 140113
rect 186801 140085 186829 140113
rect 186739 140023 186767 140051
rect 186801 140023 186829 140051
rect 186739 139961 186767 139989
rect 186801 139961 186829 139989
rect 202099 140147 202127 140175
rect 202161 140147 202189 140175
rect 202099 140085 202127 140113
rect 202161 140085 202189 140113
rect 202099 140023 202127 140051
rect 202161 140023 202189 140051
rect 202099 139961 202127 139989
rect 202161 139961 202189 139989
rect 217459 140147 217487 140175
rect 217521 140147 217549 140175
rect 217459 140085 217487 140113
rect 217521 140085 217549 140113
rect 217459 140023 217487 140051
rect 217521 140023 217549 140051
rect 217459 139961 217487 139989
rect 217521 139961 217549 139989
rect 232819 140147 232847 140175
rect 232881 140147 232909 140175
rect 232819 140085 232847 140113
rect 232881 140085 232909 140113
rect 232819 140023 232847 140051
rect 232881 140023 232909 140051
rect 232819 139961 232847 139989
rect 232881 139961 232909 139989
rect 248179 140147 248207 140175
rect 248241 140147 248269 140175
rect 248179 140085 248207 140113
rect 248241 140085 248269 140113
rect 248179 140023 248207 140051
rect 248241 140023 248269 140051
rect 248179 139961 248207 139989
rect 248241 139961 248269 139989
rect 263539 140147 263567 140175
rect 263601 140147 263629 140175
rect 263539 140085 263567 140113
rect 263601 140085 263629 140113
rect 263539 140023 263567 140051
rect 263601 140023 263629 140051
rect 263539 139961 263567 139989
rect 263601 139961 263629 139989
rect 278899 140147 278927 140175
rect 278961 140147 278989 140175
rect 278899 140085 278927 140113
rect 278961 140085 278989 140113
rect 278899 140023 278927 140051
rect 278961 140023 278989 140051
rect 278899 139961 278927 139989
rect 278961 139961 278989 139989
rect 102259 137147 102287 137175
rect 102321 137147 102349 137175
rect 102259 137085 102287 137113
rect 102321 137085 102349 137113
rect 102259 137023 102287 137051
rect 102321 137023 102349 137051
rect 102259 136961 102287 136989
rect 102321 136961 102349 136989
rect 117619 137147 117647 137175
rect 117681 137147 117709 137175
rect 117619 137085 117647 137113
rect 117681 137085 117709 137113
rect 117619 137023 117647 137051
rect 117681 137023 117709 137051
rect 117619 136961 117647 136989
rect 117681 136961 117709 136989
rect 132979 137147 133007 137175
rect 133041 137147 133069 137175
rect 132979 137085 133007 137113
rect 133041 137085 133069 137113
rect 132979 137023 133007 137051
rect 133041 137023 133069 137051
rect 132979 136961 133007 136989
rect 133041 136961 133069 136989
rect 148339 137147 148367 137175
rect 148401 137147 148429 137175
rect 148339 137085 148367 137113
rect 148401 137085 148429 137113
rect 148339 137023 148367 137051
rect 148401 137023 148429 137051
rect 148339 136961 148367 136989
rect 148401 136961 148429 136989
rect 163699 137147 163727 137175
rect 163761 137147 163789 137175
rect 163699 137085 163727 137113
rect 163761 137085 163789 137113
rect 163699 137023 163727 137051
rect 163761 137023 163789 137051
rect 163699 136961 163727 136989
rect 163761 136961 163789 136989
rect 179059 137147 179087 137175
rect 179121 137147 179149 137175
rect 179059 137085 179087 137113
rect 179121 137085 179149 137113
rect 179059 137023 179087 137051
rect 179121 137023 179149 137051
rect 179059 136961 179087 136989
rect 179121 136961 179149 136989
rect 194419 137147 194447 137175
rect 194481 137147 194509 137175
rect 194419 137085 194447 137113
rect 194481 137085 194509 137113
rect 194419 137023 194447 137051
rect 194481 137023 194509 137051
rect 194419 136961 194447 136989
rect 194481 136961 194509 136989
rect 209779 137147 209807 137175
rect 209841 137147 209869 137175
rect 209779 137085 209807 137113
rect 209841 137085 209869 137113
rect 209779 137023 209807 137051
rect 209841 137023 209869 137051
rect 209779 136961 209807 136989
rect 209841 136961 209869 136989
rect 225139 137147 225167 137175
rect 225201 137147 225229 137175
rect 225139 137085 225167 137113
rect 225201 137085 225229 137113
rect 225139 137023 225167 137051
rect 225201 137023 225229 137051
rect 225139 136961 225167 136989
rect 225201 136961 225229 136989
rect 240499 137147 240527 137175
rect 240561 137147 240589 137175
rect 240499 137085 240527 137113
rect 240561 137085 240589 137113
rect 240499 137023 240527 137051
rect 240561 137023 240589 137051
rect 240499 136961 240527 136989
rect 240561 136961 240589 136989
rect 255859 137147 255887 137175
rect 255921 137147 255949 137175
rect 255859 137085 255887 137113
rect 255921 137085 255949 137113
rect 255859 137023 255887 137051
rect 255921 137023 255949 137051
rect 255859 136961 255887 136989
rect 255921 136961 255949 136989
rect 271219 137147 271247 137175
rect 271281 137147 271309 137175
rect 271219 137085 271247 137113
rect 271281 137085 271309 137113
rect 271219 137023 271247 137051
rect 271281 137023 271309 137051
rect 271219 136961 271247 136989
rect 271281 136961 271309 136989
rect 279237 137147 279265 137175
rect 279299 137147 279327 137175
rect 279361 137147 279389 137175
rect 279423 137147 279451 137175
rect 279237 137085 279265 137113
rect 279299 137085 279327 137113
rect 279361 137085 279389 137113
rect 279423 137085 279451 137113
rect 279237 137023 279265 137051
rect 279299 137023 279327 137051
rect 279361 137023 279389 137051
rect 279423 137023 279451 137051
rect 279237 136961 279265 136989
rect 279299 136961 279327 136989
rect 279361 136961 279389 136989
rect 279423 136961 279451 136989
rect 109939 131147 109967 131175
rect 110001 131147 110029 131175
rect 109939 131085 109967 131113
rect 110001 131085 110029 131113
rect 109939 131023 109967 131051
rect 110001 131023 110029 131051
rect 109939 130961 109967 130989
rect 110001 130961 110029 130989
rect 125299 131147 125327 131175
rect 125361 131147 125389 131175
rect 125299 131085 125327 131113
rect 125361 131085 125389 131113
rect 125299 131023 125327 131051
rect 125361 131023 125389 131051
rect 125299 130961 125327 130989
rect 125361 130961 125389 130989
rect 140659 131147 140687 131175
rect 140721 131147 140749 131175
rect 140659 131085 140687 131113
rect 140721 131085 140749 131113
rect 140659 131023 140687 131051
rect 140721 131023 140749 131051
rect 140659 130961 140687 130989
rect 140721 130961 140749 130989
rect 156019 131147 156047 131175
rect 156081 131147 156109 131175
rect 156019 131085 156047 131113
rect 156081 131085 156109 131113
rect 156019 131023 156047 131051
rect 156081 131023 156109 131051
rect 156019 130961 156047 130989
rect 156081 130961 156109 130989
rect 171379 131147 171407 131175
rect 171441 131147 171469 131175
rect 171379 131085 171407 131113
rect 171441 131085 171469 131113
rect 171379 131023 171407 131051
rect 171441 131023 171469 131051
rect 171379 130961 171407 130989
rect 171441 130961 171469 130989
rect 186739 131147 186767 131175
rect 186801 131147 186829 131175
rect 186739 131085 186767 131113
rect 186801 131085 186829 131113
rect 186739 131023 186767 131051
rect 186801 131023 186829 131051
rect 186739 130961 186767 130989
rect 186801 130961 186829 130989
rect 202099 131147 202127 131175
rect 202161 131147 202189 131175
rect 202099 131085 202127 131113
rect 202161 131085 202189 131113
rect 202099 131023 202127 131051
rect 202161 131023 202189 131051
rect 202099 130961 202127 130989
rect 202161 130961 202189 130989
rect 217459 131147 217487 131175
rect 217521 131147 217549 131175
rect 217459 131085 217487 131113
rect 217521 131085 217549 131113
rect 217459 131023 217487 131051
rect 217521 131023 217549 131051
rect 217459 130961 217487 130989
rect 217521 130961 217549 130989
rect 232819 131147 232847 131175
rect 232881 131147 232909 131175
rect 232819 131085 232847 131113
rect 232881 131085 232909 131113
rect 232819 131023 232847 131051
rect 232881 131023 232909 131051
rect 232819 130961 232847 130989
rect 232881 130961 232909 130989
rect 248179 131147 248207 131175
rect 248241 131147 248269 131175
rect 248179 131085 248207 131113
rect 248241 131085 248269 131113
rect 248179 131023 248207 131051
rect 248241 131023 248269 131051
rect 248179 130961 248207 130989
rect 248241 130961 248269 130989
rect 263539 131147 263567 131175
rect 263601 131147 263629 131175
rect 263539 131085 263567 131113
rect 263601 131085 263629 131113
rect 263539 131023 263567 131051
rect 263601 131023 263629 131051
rect 263539 130961 263567 130989
rect 263601 130961 263629 130989
rect 278899 131147 278927 131175
rect 278961 131147 278989 131175
rect 278899 131085 278927 131113
rect 278961 131085 278989 131113
rect 278899 131023 278927 131051
rect 278961 131023 278989 131051
rect 278899 130961 278927 130989
rect 278961 130961 278989 130989
rect 102259 128147 102287 128175
rect 102321 128147 102349 128175
rect 102259 128085 102287 128113
rect 102321 128085 102349 128113
rect 102259 128023 102287 128051
rect 102321 128023 102349 128051
rect 102259 127961 102287 127989
rect 102321 127961 102349 127989
rect 117619 128147 117647 128175
rect 117681 128147 117709 128175
rect 117619 128085 117647 128113
rect 117681 128085 117709 128113
rect 117619 128023 117647 128051
rect 117681 128023 117709 128051
rect 117619 127961 117647 127989
rect 117681 127961 117709 127989
rect 132979 128147 133007 128175
rect 133041 128147 133069 128175
rect 132979 128085 133007 128113
rect 133041 128085 133069 128113
rect 132979 128023 133007 128051
rect 133041 128023 133069 128051
rect 132979 127961 133007 127989
rect 133041 127961 133069 127989
rect 148339 128147 148367 128175
rect 148401 128147 148429 128175
rect 148339 128085 148367 128113
rect 148401 128085 148429 128113
rect 148339 128023 148367 128051
rect 148401 128023 148429 128051
rect 148339 127961 148367 127989
rect 148401 127961 148429 127989
rect 163699 128147 163727 128175
rect 163761 128147 163789 128175
rect 163699 128085 163727 128113
rect 163761 128085 163789 128113
rect 163699 128023 163727 128051
rect 163761 128023 163789 128051
rect 163699 127961 163727 127989
rect 163761 127961 163789 127989
rect 179059 128147 179087 128175
rect 179121 128147 179149 128175
rect 179059 128085 179087 128113
rect 179121 128085 179149 128113
rect 179059 128023 179087 128051
rect 179121 128023 179149 128051
rect 179059 127961 179087 127989
rect 179121 127961 179149 127989
rect 194419 128147 194447 128175
rect 194481 128147 194509 128175
rect 194419 128085 194447 128113
rect 194481 128085 194509 128113
rect 194419 128023 194447 128051
rect 194481 128023 194509 128051
rect 194419 127961 194447 127989
rect 194481 127961 194509 127989
rect 209779 128147 209807 128175
rect 209841 128147 209869 128175
rect 209779 128085 209807 128113
rect 209841 128085 209869 128113
rect 209779 128023 209807 128051
rect 209841 128023 209869 128051
rect 209779 127961 209807 127989
rect 209841 127961 209869 127989
rect 225139 128147 225167 128175
rect 225201 128147 225229 128175
rect 225139 128085 225167 128113
rect 225201 128085 225229 128113
rect 225139 128023 225167 128051
rect 225201 128023 225229 128051
rect 225139 127961 225167 127989
rect 225201 127961 225229 127989
rect 240499 128147 240527 128175
rect 240561 128147 240589 128175
rect 240499 128085 240527 128113
rect 240561 128085 240589 128113
rect 240499 128023 240527 128051
rect 240561 128023 240589 128051
rect 240499 127961 240527 127989
rect 240561 127961 240589 127989
rect 255859 128147 255887 128175
rect 255921 128147 255949 128175
rect 255859 128085 255887 128113
rect 255921 128085 255949 128113
rect 255859 128023 255887 128051
rect 255921 128023 255949 128051
rect 255859 127961 255887 127989
rect 255921 127961 255949 127989
rect 271219 128147 271247 128175
rect 271281 128147 271309 128175
rect 271219 128085 271247 128113
rect 271281 128085 271309 128113
rect 271219 128023 271247 128051
rect 271281 128023 271309 128051
rect 271219 127961 271247 127989
rect 271281 127961 271309 127989
rect 279237 128147 279265 128175
rect 279299 128147 279327 128175
rect 279361 128147 279389 128175
rect 279423 128147 279451 128175
rect 279237 128085 279265 128113
rect 279299 128085 279327 128113
rect 279361 128085 279389 128113
rect 279423 128085 279451 128113
rect 279237 128023 279265 128051
rect 279299 128023 279327 128051
rect 279361 128023 279389 128051
rect 279423 128023 279451 128051
rect 279237 127961 279265 127989
rect 279299 127961 279327 127989
rect 279361 127961 279389 127989
rect 279423 127961 279451 127989
rect 109939 122147 109967 122175
rect 110001 122147 110029 122175
rect 109939 122085 109967 122113
rect 110001 122085 110029 122113
rect 109939 122023 109967 122051
rect 110001 122023 110029 122051
rect 109939 121961 109967 121989
rect 110001 121961 110029 121989
rect 125299 122147 125327 122175
rect 125361 122147 125389 122175
rect 125299 122085 125327 122113
rect 125361 122085 125389 122113
rect 125299 122023 125327 122051
rect 125361 122023 125389 122051
rect 125299 121961 125327 121989
rect 125361 121961 125389 121989
rect 140659 122147 140687 122175
rect 140721 122147 140749 122175
rect 140659 122085 140687 122113
rect 140721 122085 140749 122113
rect 140659 122023 140687 122051
rect 140721 122023 140749 122051
rect 140659 121961 140687 121989
rect 140721 121961 140749 121989
rect 156019 122147 156047 122175
rect 156081 122147 156109 122175
rect 156019 122085 156047 122113
rect 156081 122085 156109 122113
rect 156019 122023 156047 122051
rect 156081 122023 156109 122051
rect 156019 121961 156047 121989
rect 156081 121961 156109 121989
rect 171379 122147 171407 122175
rect 171441 122147 171469 122175
rect 171379 122085 171407 122113
rect 171441 122085 171469 122113
rect 171379 122023 171407 122051
rect 171441 122023 171469 122051
rect 171379 121961 171407 121989
rect 171441 121961 171469 121989
rect 186739 122147 186767 122175
rect 186801 122147 186829 122175
rect 186739 122085 186767 122113
rect 186801 122085 186829 122113
rect 186739 122023 186767 122051
rect 186801 122023 186829 122051
rect 186739 121961 186767 121989
rect 186801 121961 186829 121989
rect 202099 122147 202127 122175
rect 202161 122147 202189 122175
rect 202099 122085 202127 122113
rect 202161 122085 202189 122113
rect 202099 122023 202127 122051
rect 202161 122023 202189 122051
rect 202099 121961 202127 121989
rect 202161 121961 202189 121989
rect 217459 122147 217487 122175
rect 217521 122147 217549 122175
rect 217459 122085 217487 122113
rect 217521 122085 217549 122113
rect 217459 122023 217487 122051
rect 217521 122023 217549 122051
rect 217459 121961 217487 121989
rect 217521 121961 217549 121989
rect 232819 122147 232847 122175
rect 232881 122147 232909 122175
rect 232819 122085 232847 122113
rect 232881 122085 232909 122113
rect 232819 122023 232847 122051
rect 232881 122023 232909 122051
rect 232819 121961 232847 121989
rect 232881 121961 232909 121989
rect 248179 122147 248207 122175
rect 248241 122147 248269 122175
rect 248179 122085 248207 122113
rect 248241 122085 248269 122113
rect 248179 122023 248207 122051
rect 248241 122023 248269 122051
rect 248179 121961 248207 121989
rect 248241 121961 248269 121989
rect 263539 122147 263567 122175
rect 263601 122147 263629 122175
rect 263539 122085 263567 122113
rect 263601 122085 263629 122113
rect 263539 122023 263567 122051
rect 263601 122023 263629 122051
rect 263539 121961 263567 121989
rect 263601 121961 263629 121989
rect 278899 122147 278927 122175
rect 278961 122147 278989 122175
rect 278899 122085 278927 122113
rect 278961 122085 278989 122113
rect 278899 122023 278927 122051
rect 278961 122023 278989 122051
rect 278899 121961 278927 121989
rect 278961 121961 278989 121989
rect 102259 119147 102287 119175
rect 102321 119147 102349 119175
rect 102259 119085 102287 119113
rect 102321 119085 102349 119113
rect 102259 119023 102287 119051
rect 102321 119023 102349 119051
rect 102259 118961 102287 118989
rect 102321 118961 102349 118989
rect 117619 119147 117647 119175
rect 117681 119147 117709 119175
rect 117619 119085 117647 119113
rect 117681 119085 117709 119113
rect 117619 119023 117647 119051
rect 117681 119023 117709 119051
rect 117619 118961 117647 118989
rect 117681 118961 117709 118989
rect 132979 119147 133007 119175
rect 133041 119147 133069 119175
rect 132979 119085 133007 119113
rect 133041 119085 133069 119113
rect 132979 119023 133007 119051
rect 133041 119023 133069 119051
rect 132979 118961 133007 118989
rect 133041 118961 133069 118989
rect 148339 119147 148367 119175
rect 148401 119147 148429 119175
rect 148339 119085 148367 119113
rect 148401 119085 148429 119113
rect 148339 119023 148367 119051
rect 148401 119023 148429 119051
rect 148339 118961 148367 118989
rect 148401 118961 148429 118989
rect 163699 119147 163727 119175
rect 163761 119147 163789 119175
rect 163699 119085 163727 119113
rect 163761 119085 163789 119113
rect 163699 119023 163727 119051
rect 163761 119023 163789 119051
rect 163699 118961 163727 118989
rect 163761 118961 163789 118989
rect 179059 119147 179087 119175
rect 179121 119147 179149 119175
rect 179059 119085 179087 119113
rect 179121 119085 179149 119113
rect 179059 119023 179087 119051
rect 179121 119023 179149 119051
rect 179059 118961 179087 118989
rect 179121 118961 179149 118989
rect 194419 119147 194447 119175
rect 194481 119147 194509 119175
rect 194419 119085 194447 119113
rect 194481 119085 194509 119113
rect 194419 119023 194447 119051
rect 194481 119023 194509 119051
rect 194419 118961 194447 118989
rect 194481 118961 194509 118989
rect 209779 119147 209807 119175
rect 209841 119147 209869 119175
rect 209779 119085 209807 119113
rect 209841 119085 209869 119113
rect 209779 119023 209807 119051
rect 209841 119023 209869 119051
rect 209779 118961 209807 118989
rect 209841 118961 209869 118989
rect 225139 119147 225167 119175
rect 225201 119147 225229 119175
rect 225139 119085 225167 119113
rect 225201 119085 225229 119113
rect 225139 119023 225167 119051
rect 225201 119023 225229 119051
rect 225139 118961 225167 118989
rect 225201 118961 225229 118989
rect 240499 119147 240527 119175
rect 240561 119147 240589 119175
rect 240499 119085 240527 119113
rect 240561 119085 240589 119113
rect 240499 119023 240527 119051
rect 240561 119023 240589 119051
rect 240499 118961 240527 118989
rect 240561 118961 240589 118989
rect 255859 119147 255887 119175
rect 255921 119147 255949 119175
rect 255859 119085 255887 119113
rect 255921 119085 255949 119113
rect 255859 119023 255887 119051
rect 255921 119023 255949 119051
rect 255859 118961 255887 118989
rect 255921 118961 255949 118989
rect 271219 119147 271247 119175
rect 271281 119147 271309 119175
rect 271219 119085 271247 119113
rect 271281 119085 271309 119113
rect 271219 119023 271247 119051
rect 271281 119023 271309 119051
rect 271219 118961 271247 118989
rect 271281 118961 271309 118989
rect 279237 119147 279265 119175
rect 279299 119147 279327 119175
rect 279361 119147 279389 119175
rect 279423 119147 279451 119175
rect 279237 119085 279265 119113
rect 279299 119085 279327 119113
rect 279361 119085 279389 119113
rect 279423 119085 279451 119113
rect 279237 119023 279265 119051
rect 279299 119023 279327 119051
rect 279361 119023 279389 119051
rect 279423 119023 279451 119051
rect 279237 118961 279265 118989
rect 279299 118961 279327 118989
rect 279361 118961 279389 118989
rect 279423 118961 279451 118989
rect 109939 113147 109967 113175
rect 110001 113147 110029 113175
rect 109939 113085 109967 113113
rect 110001 113085 110029 113113
rect 109939 113023 109967 113051
rect 110001 113023 110029 113051
rect 109939 112961 109967 112989
rect 110001 112961 110029 112989
rect 125299 113147 125327 113175
rect 125361 113147 125389 113175
rect 125299 113085 125327 113113
rect 125361 113085 125389 113113
rect 125299 113023 125327 113051
rect 125361 113023 125389 113051
rect 125299 112961 125327 112989
rect 125361 112961 125389 112989
rect 140659 113147 140687 113175
rect 140721 113147 140749 113175
rect 140659 113085 140687 113113
rect 140721 113085 140749 113113
rect 140659 113023 140687 113051
rect 140721 113023 140749 113051
rect 140659 112961 140687 112989
rect 140721 112961 140749 112989
rect 156019 113147 156047 113175
rect 156081 113147 156109 113175
rect 156019 113085 156047 113113
rect 156081 113085 156109 113113
rect 156019 113023 156047 113051
rect 156081 113023 156109 113051
rect 156019 112961 156047 112989
rect 156081 112961 156109 112989
rect 171379 113147 171407 113175
rect 171441 113147 171469 113175
rect 171379 113085 171407 113113
rect 171441 113085 171469 113113
rect 171379 113023 171407 113051
rect 171441 113023 171469 113051
rect 171379 112961 171407 112989
rect 171441 112961 171469 112989
rect 186739 113147 186767 113175
rect 186801 113147 186829 113175
rect 186739 113085 186767 113113
rect 186801 113085 186829 113113
rect 186739 113023 186767 113051
rect 186801 113023 186829 113051
rect 186739 112961 186767 112989
rect 186801 112961 186829 112989
rect 202099 113147 202127 113175
rect 202161 113147 202189 113175
rect 202099 113085 202127 113113
rect 202161 113085 202189 113113
rect 202099 113023 202127 113051
rect 202161 113023 202189 113051
rect 202099 112961 202127 112989
rect 202161 112961 202189 112989
rect 217459 113147 217487 113175
rect 217521 113147 217549 113175
rect 217459 113085 217487 113113
rect 217521 113085 217549 113113
rect 217459 113023 217487 113051
rect 217521 113023 217549 113051
rect 217459 112961 217487 112989
rect 217521 112961 217549 112989
rect 232819 113147 232847 113175
rect 232881 113147 232909 113175
rect 232819 113085 232847 113113
rect 232881 113085 232909 113113
rect 232819 113023 232847 113051
rect 232881 113023 232909 113051
rect 232819 112961 232847 112989
rect 232881 112961 232909 112989
rect 248179 113147 248207 113175
rect 248241 113147 248269 113175
rect 248179 113085 248207 113113
rect 248241 113085 248269 113113
rect 248179 113023 248207 113051
rect 248241 113023 248269 113051
rect 248179 112961 248207 112989
rect 248241 112961 248269 112989
rect 263539 113147 263567 113175
rect 263601 113147 263629 113175
rect 263539 113085 263567 113113
rect 263601 113085 263629 113113
rect 263539 113023 263567 113051
rect 263601 113023 263629 113051
rect 263539 112961 263567 112989
rect 263601 112961 263629 112989
rect 278899 113147 278927 113175
rect 278961 113147 278989 113175
rect 278899 113085 278927 113113
rect 278961 113085 278989 113113
rect 278899 113023 278927 113051
rect 278961 113023 278989 113051
rect 278899 112961 278927 112989
rect 278961 112961 278989 112989
rect 102259 110147 102287 110175
rect 102321 110147 102349 110175
rect 102259 110085 102287 110113
rect 102321 110085 102349 110113
rect 102259 110023 102287 110051
rect 102321 110023 102349 110051
rect 102259 109961 102287 109989
rect 102321 109961 102349 109989
rect 117619 110147 117647 110175
rect 117681 110147 117709 110175
rect 117619 110085 117647 110113
rect 117681 110085 117709 110113
rect 117619 110023 117647 110051
rect 117681 110023 117709 110051
rect 117619 109961 117647 109989
rect 117681 109961 117709 109989
rect 132979 110147 133007 110175
rect 133041 110147 133069 110175
rect 132979 110085 133007 110113
rect 133041 110085 133069 110113
rect 132979 110023 133007 110051
rect 133041 110023 133069 110051
rect 132979 109961 133007 109989
rect 133041 109961 133069 109989
rect 148339 110147 148367 110175
rect 148401 110147 148429 110175
rect 148339 110085 148367 110113
rect 148401 110085 148429 110113
rect 148339 110023 148367 110051
rect 148401 110023 148429 110051
rect 148339 109961 148367 109989
rect 148401 109961 148429 109989
rect 163699 110147 163727 110175
rect 163761 110147 163789 110175
rect 163699 110085 163727 110113
rect 163761 110085 163789 110113
rect 163699 110023 163727 110051
rect 163761 110023 163789 110051
rect 163699 109961 163727 109989
rect 163761 109961 163789 109989
rect 179059 110147 179087 110175
rect 179121 110147 179149 110175
rect 179059 110085 179087 110113
rect 179121 110085 179149 110113
rect 179059 110023 179087 110051
rect 179121 110023 179149 110051
rect 179059 109961 179087 109989
rect 179121 109961 179149 109989
rect 194419 110147 194447 110175
rect 194481 110147 194509 110175
rect 194419 110085 194447 110113
rect 194481 110085 194509 110113
rect 194419 110023 194447 110051
rect 194481 110023 194509 110051
rect 194419 109961 194447 109989
rect 194481 109961 194509 109989
rect 209779 110147 209807 110175
rect 209841 110147 209869 110175
rect 209779 110085 209807 110113
rect 209841 110085 209869 110113
rect 209779 110023 209807 110051
rect 209841 110023 209869 110051
rect 209779 109961 209807 109989
rect 209841 109961 209869 109989
rect 225139 110147 225167 110175
rect 225201 110147 225229 110175
rect 225139 110085 225167 110113
rect 225201 110085 225229 110113
rect 225139 110023 225167 110051
rect 225201 110023 225229 110051
rect 225139 109961 225167 109989
rect 225201 109961 225229 109989
rect 240499 110147 240527 110175
rect 240561 110147 240589 110175
rect 240499 110085 240527 110113
rect 240561 110085 240589 110113
rect 240499 110023 240527 110051
rect 240561 110023 240589 110051
rect 240499 109961 240527 109989
rect 240561 109961 240589 109989
rect 255859 110147 255887 110175
rect 255921 110147 255949 110175
rect 255859 110085 255887 110113
rect 255921 110085 255949 110113
rect 255859 110023 255887 110051
rect 255921 110023 255949 110051
rect 255859 109961 255887 109989
rect 255921 109961 255949 109989
rect 271219 110147 271247 110175
rect 271281 110147 271309 110175
rect 271219 110085 271247 110113
rect 271281 110085 271309 110113
rect 271219 110023 271247 110051
rect 271281 110023 271309 110051
rect 271219 109961 271247 109989
rect 271281 109961 271309 109989
rect 279237 110147 279265 110175
rect 279299 110147 279327 110175
rect 279361 110147 279389 110175
rect 279423 110147 279451 110175
rect 279237 110085 279265 110113
rect 279299 110085 279327 110113
rect 279361 110085 279389 110113
rect 279423 110085 279451 110113
rect 279237 110023 279265 110051
rect 279299 110023 279327 110051
rect 279361 110023 279389 110051
rect 279423 110023 279451 110051
rect 279237 109961 279265 109989
rect 279299 109961 279327 109989
rect 279361 109961 279389 109989
rect 279423 109961 279451 109989
rect 109939 104147 109967 104175
rect 110001 104147 110029 104175
rect 109939 104085 109967 104113
rect 110001 104085 110029 104113
rect 109939 104023 109967 104051
rect 110001 104023 110029 104051
rect 109939 103961 109967 103989
rect 110001 103961 110029 103989
rect 125299 104147 125327 104175
rect 125361 104147 125389 104175
rect 125299 104085 125327 104113
rect 125361 104085 125389 104113
rect 125299 104023 125327 104051
rect 125361 104023 125389 104051
rect 125299 103961 125327 103989
rect 125361 103961 125389 103989
rect 140659 104147 140687 104175
rect 140721 104147 140749 104175
rect 140659 104085 140687 104113
rect 140721 104085 140749 104113
rect 140659 104023 140687 104051
rect 140721 104023 140749 104051
rect 140659 103961 140687 103989
rect 140721 103961 140749 103989
rect 156019 104147 156047 104175
rect 156081 104147 156109 104175
rect 156019 104085 156047 104113
rect 156081 104085 156109 104113
rect 156019 104023 156047 104051
rect 156081 104023 156109 104051
rect 156019 103961 156047 103989
rect 156081 103961 156109 103989
rect 171379 104147 171407 104175
rect 171441 104147 171469 104175
rect 171379 104085 171407 104113
rect 171441 104085 171469 104113
rect 171379 104023 171407 104051
rect 171441 104023 171469 104051
rect 171379 103961 171407 103989
rect 171441 103961 171469 103989
rect 186739 104147 186767 104175
rect 186801 104147 186829 104175
rect 186739 104085 186767 104113
rect 186801 104085 186829 104113
rect 186739 104023 186767 104051
rect 186801 104023 186829 104051
rect 186739 103961 186767 103989
rect 186801 103961 186829 103989
rect 202099 104147 202127 104175
rect 202161 104147 202189 104175
rect 202099 104085 202127 104113
rect 202161 104085 202189 104113
rect 202099 104023 202127 104051
rect 202161 104023 202189 104051
rect 202099 103961 202127 103989
rect 202161 103961 202189 103989
rect 217459 104147 217487 104175
rect 217521 104147 217549 104175
rect 217459 104085 217487 104113
rect 217521 104085 217549 104113
rect 217459 104023 217487 104051
rect 217521 104023 217549 104051
rect 217459 103961 217487 103989
rect 217521 103961 217549 103989
rect 232819 104147 232847 104175
rect 232881 104147 232909 104175
rect 232819 104085 232847 104113
rect 232881 104085 232909 104113
rect 232819 104023 232847 104051
rect 232881 104023 232909 104051
rect 232819 103961 232847 103989
rect 232881 103961 232909 103989
rect 248179 104147 248207 104175
rect 248241 104147 248269 104175
rect 248179 104085 248207 104113
rect 248241 104085 248269 104113
rect 248179 104023 248207 104051
rect 248241 104023 248269 104051
rect 248179 103961 248207 103989
rect 248241 103961 248269 103989
rect 263539 104147 263567 104175
rect 263601 104147 263629 104175
rect 263539 104085 263567 104113
rect 263601 104085 263629 104113
rect 263539 104023 263567 104051
rect 263601 104023 263629 104051
rect 263539 103961 263567 103989
rect 263601 103961 263629 103989
rect 278899 104147 278927 104175
rect 278961 104147 278989 104175
rect 278899 104085 278927 104113
rect 278961 104085 278989 104113
rect 278899 104023 278927 104051
rect 278961 104023 278989 104051
rect 278899 103961 278927 103989
rect 278961 103961 278989 103989
rect 279237 101147 279265 101175
rect 279299 101147 279327 101175
rect 279361 101147 279389 101175
rect 279423 101147 279451 101175
rect 279237 101085 279265 101113
rect 279299 101085 279327 101113
rect 279361 101085 279389 101113
rect 279423 101085 279451 101113
rect 279237 101023 279265 101051
rect 279299 101023 279327 101051
rect 279361 101023 279389 101051
rect 279423 101023 279451 101051
rect 279237 100961 279265 100989
rect 279299 100961 279327 100989
rect 279361 100961 279389 100989
rect 279423 100961 279451 100989
rect 110277 92147 110305 92175
rect 110339 92147 110367 92175
rect 110401 92147 110429 92175
rect 110463 92147 110491 92175
rect 110277 92085 110305 92113
rect 110339 92085 110367 92113
rect 110401 92085 110429 92113
rect 110463 92085 110491 92113
rect 110277 92023 110305 92051
rect 110339 92023 110367 92051
rect 110401 92023 110429 92051
rect 110463 92023 110491 92051
rect 110277 91961 110305 91989
rect 110339 91961 110367 91989
rect 110401 91961 110429 91989
rect 110463 91961 110491 91989
rect 110277 83147 110305 83175
rect 110339 83147 110367 83175
rect 110401 83147 110429 83175
rect 110463 83147 110491 83175
rect 110277 83085 110305 83113
rect 110339 83085 110367 83113
rect 110401 83085 110429 83113
rect 110463 83085 110491 83113
rect 110277 83023 110305 83051
rect 110339 83023 110367 83051
rect 110401 83023 110429 83051
rect 110463 83023 110491 83051
rect 110277 82961 110305 82989
rect 110339 82961 110367 82989
rect 110401 82961 110429 82989
rect 110463 82961 110491 82989
rect 110277 74147 110305 74175
rect 110339 74147 110367 74175
rect 110401 74147 110429 74175
rect 110463 74147 110491 74175
rect 110277 74085 110305 74113
rect 110339 74085 110367 74113
rect 110401 74085 110429 74113
rect 110463 74085 110491 74113
rect 110277 74023 110305 74051
rect 110339 74023 110367 74051
rect 110401 74023 110429 74051
rect 110463 74023 110491 74051
rect 110277 73961 110305 73989
rect 110339 73961 110367 73989
rect 110401 73961 110429 73989
rect 110463 73961 110491 73989
rect 110277 65147 110305 65175
rect 110339 65147 110367 65175
rect 110401 65147 110429 65175
rect 110463 65147 110491 65175
rect 110277 65085 110305 65113
rect 110339 65085 110367 65113
rect 110401 65085 110429 65113
rect 110463 65085 110491 65113
rect 110277 65023 110305 65051
rect 110339 65023 110367 65051
rect 110401 65023 110429 65051
rect 110463 65023 110491 65051
rect 110277 64961 110305 64989
rect 110339 64961 110367 64989
rect 110401 64961 110429 64989
rect 110463 64961 110491 64989
rect 110277 56147 110305 56175
rect 110339 56147 110367 56175
rect 110401 56147 110429 56175
rect 110463 56147 110491 56175
rect 110277 56085 110305 56113
rect 110339 56085 110367 56113
rect 110401 56085 110429 56113
rect 110463 56085 110491 56113
rect 110277 56023 110305 56051
rect 110339 56023 110367 56051
rect 110401 56023 110429 56051
rect 110463 56023 110491 56051
rect 110277 55961 110305 55989
rect 110339 55961 110367 55989
rect 110401 55961 110429 55989
rect 110463 55961 110491 55989
rect 110277 47147 110305 47175
rect 110339 47147 110367 47175
rect 110401 47147 110429 47175
rect 110463 47147 110491 47175
rect 110277 47085 110305 47113
rect 110339 47085 110367 47113
rect 110401 47085 110429 47113
rect 110463 47085 110491 47113
rect 110277 47023 110305 47051
rect 110339 47023 110367 47051
rect 110401 47023 110429 47051
rect 110463 47023 110491 47051
rect 110277 46961 110305 46989
rect 110339 46961 110367 46989
rect 110401 46961 110429 46989
rect 110463 46961 110491 46989
rect 110277 38147 110305 38175
rect 110339 38147 110367 38175
rect 110401 38147 110429 38175
rect 110463 38147 110491 38175
rect 110277 38085 110305 38113
rect 110339 38085 110367 38113
rect 110401 38085 110429 38113
rect 110463 38085 110491 38113
rect 110277 38023 110305 38051
rect 110339 38023 110367 38051
rect 110401 38023 110429 38051
rect 110463 38023 110491 38051
rect 110277 37961 110305 37989
rect 110339 37961 110367 37989
rect 110401 37961 110429 37989
rect 110463 37961 110491 37989
rect 110277 29147 110305 29175
rect 110339 29147 110367 29175
rect 110401 29147 110429 29175
rect 110463 29147 110491 29175
rect 110277 29085 110305 29113
rect 110339 29085 110367 29113
rect 110401 29085 110429 29113
rect 110463 29085 110491 29113
rect 110277 29023 110305 29051
rect 110339 29023 110367 29051
rect 110401 29023 110429 29051
rect 110463 29023 110491 29051
rect 110277 28961 110305 28989
rect 110339 28961 110367 28989
rect 110401 28961 110429 28989
rect 110463 28961 110491 28989
rect 110277 20147 110305 20175
rect 110339 20147 110367 20175
rect 110401 20147 110429 20175
rect 110463 20147 110491 20175
rect 110277 20085 110305 20113
rect 110339 20085 110367 20113
rect 110401 20085 110429 20113
rect 110463 20085 110491 20113
rect 110277 20023 110305 20051
rect 110339 20023 110367 20051
rect 110401 20023 110429 20051
rect 110463 20023 110491 20051
rect 110277 19961 110305 19989
rect 110339 19961 110367 19989
rect 110401 19961 110429 19989
rect 110463 19961 110491 19989
rect 96777 14147 96805 14175
rect 96839 14147 96867 14175
rect 96901 14147 96929 14175
rect 96963 14147 96991 14175
rect 96777 14085 96805 14113
rect 96839 14085 96867 14113
rect 96901 14085 96929 14113
rect 96963 14085 96991 14113
rect 96777 14023 96805 14051
rect 96839 14023 96867 14051
rect 96901 14023 96929 14051
rect 96963 14023 96991 14051
rect 96777 13961 96805 13989
rect 96839 13961 96867 13989
rect 96901 13961 96929 13989
rect 96963 13961 96991 13989
rect 96777 5147 96805 5175
rect 96839 5147 96867 5175
rect 96901 5147 96929 5175
rect 96963 5147 96991 5175
rect 96777 5085 96805 5113
rect 96839 5085 96867 5113
rect 96901 5085 96929 5113
rect 96963 5085 96991 5113
rect 96777 5023 96805 5051
rect 96839 5023 96867 5051
rect 96901 5023 96929 5051
rect 96963 5023 96991 5051
rect 96777 4961 96805 4989
rect 96839 4961 96867 4989
rect 96901 4961 96929 4989
rect 96963 4961 96991 4989
rect 96777 -588 96805 -560
rect 96839 -588 96867 -560
rect 96901 -588 96929 -560
rect 96963 -588 96991 -560
rect 96777 -650 96805 -622
rect 96839 -650 96867 -622
rect 96901 -650 96929 -622
rect 96963 -650 96991 -622
rect 96777 -712 96805 -684
rect 96839 -712 96867 -684
rect 96901 -712 96929 -684
rect 96963 -712 96991 -684
rect 96777 -774 96805 -746
rect 96839 -774 96867 -746
rect 96901 -774 96929 -746
rect 96963 -774 96991 -746
rect 110277 11147 110305 11175
rect 110339 11147 110367 11175
rect 110401 11147 110429 11175
rect 110463 11147 110491 11175
rect 110277 11085 110305 11113
rect 110339 11085 110367 11113
rect 110401 11085 110429 11113
rect 110463 11085 110491 11113
rect 110277 11023 110305 11051
rect 110339 11023 110367 11051
rect 110401 11023 110429 11051
rect 110463 11023 110491 11051
rect 110277 10961 110305 10989
rect 110339 10961 110367 10989
rect 110401 10961 110429 10989
rect 110463 10961 110491 10989
rect 110277 2147 110305 2175
rect 110339 2147 110367 2175
rect 110401 2147 110429 2175
rect 110463 2147 110491 2175
rect 110277 2085 110305 2113
rect 110339 2085 110367 2113
rect 110401 2085 110429 2113
rect 110463 2085 110491 2113
rect 110277 2023 110305 2051
rect 110339 2023 110367 2051
rect 110401 2023 110429 2051
rect 110463 2023 110491 2051
rect 110277 1961 110305 1989
rect 110339 1961 110367 1989
rect 110401 1961 110429 1989
rect 110463 1961 110491 1989
rect 110277 -108 110305 -80
rect 110339 -108 110367 -80
rect 110401 -108 110429 -80
rect 110463 -108 110491 -80
rect 110277 -170 110305 -142
rect 110339 -170 110367 -142
rect 110401 -170 110429 -142
rect 110463 -170 110491 -142
rect 110277 -232 110305 -204
rect 110339 -232 110367 -204
rect 110401 -232 110429 -204
rect 110463 -232 110491 -204
rect 110277 -294 110305 -266
rect 110339 -294 110367 -266
rect 110401 -294 110429 -266
rect 110463 -294 110491 -266
rect 112137 95147 112165 95175
rect 112199 95147 112227 95175
rect 112261 95147 112289 95175
rect 112323 95147 112351 95175
rect 112137 95085 112165 95113
rect 112199 95085 112227 95113
rect 112261 95085 112289 95113
rect 112323 95085 112351 95113
rect 112137 95023 112165 95051
rect 112199 95023 112227 95051
rect 112261 95023 112289 95051
rect 112323 95023 112351 95051
rect 112137 94961 112165 94989
rect 112199 94961 112227 94989
rect 112261 94961 112289 94989
rect 112323 94961 112351 94989
rect 112137 86147 112165 86175
rect 112199 86147 112227 86175
rect 112261 86147 112289 86175
rect 112323 86147 112351 86175
rect 112137 86085 112165 86113
rect 112199 86085 112227 86113
rect 112261 86085 112289 86113
rect 112323 86085 112351 86113
rect 112137 86023 112165 86051
rect 112199 86023 112227 86051
rect 112261 86023 112289 86051
rect 112323 86023 112351 86051
rect 112137 85961 112165 85989
rect 112199 85961 112227 85989
rect 112261 85961 112289 85989
rect 112323 85961 112351 85989
rect 112137 77147 112165 77175
rect 112199 77147 112227 77175
rect 112261 77147 112289 77175
rect 112323 77147 112351 77175
rect 112137 77085 112165 77113
rect 112199 77085 112227 77113
rect 112261 77085 112289 77113
rect 112323 77085 112351 77113
rect 112137 77023 112165 77051
rect 112199 77023 112227 77051
rect 112261 77023 112289 77051
rect 112323 77023 112351 77051
rect 112137 76961 112165 76989
rect 112199 76961 112227 76989
rect 112261 76961 112289 76989
rect 112323 76961 112351 76989
rect 112137 68147 112165 68175
rect 112199 68147 112227 68175
rect 112261 68147 112289 68175
rect 112323 68147 112351 68175
rect 112137 68085 112165 68113
rect 112199 68085 112227 68113
rect 112261 68085 112289 68113
rect 112323 68085 112351 68113
rect 112137 68023 112165 68051
rect 112199 68023 112227 68051
rect 112261 68023 112289 68051
rect 112323 68023 112351 68051
rect 112137 67961 112165 67989
rect 112199 67961 112227 67989
rect 112261 67961 112289 67989
rect 112323 67961 112351 67989
rect 112137 59147 112165 59175
rect 112199 59147 112227 59175
rect 112261 59147 112289 59175
rect 112323 59147 112351 59175
rect 112137 59085 112165 59113
rect 112199 59085 112227 59113
rect 112261 59085 112289 59113
rect 112323 59085 112351 59113
rect 112137 59023 112165 59051
rect 112199 59023 112227 59051
rect 112261 59023 112289 59051
rect 112323 59023 112351 59051
rect 112137 58961 112165 58989
rect 112199 58961 112227 58989
rect 112261 58961 112289 58989
rect 112323 58961 112351 58989
rect 112137 50147 112165 50175
rect 112199 50147 112227 50175
rect 112261 50147 112289 50175
rect 112323 50147 112351 50175
rect 112137 50085 112165 50113
rect 112199 50085 112227 50113
rect 112261 50085 112289 50113
rect 112323 50085 112351 50113
rect 112137 50023 112165 50051
rect 112199 50023 112227 50051
rect 112261 50023 112289 50051
rect 112323 50023 112351 50051
rect 112137 49961 112165 49989
rect 112199 49961 112227 49989
rect 112261 49961 112289 49989
rect 112323 49961 112351 49989
rect 112137 41147 112165 41175
rect 112199 41147 112227 41175
rect 112261 41147 112289 41175
rect 112323 41147 112351 41175
rect 112137 41085 112165 41113
rect 112199 41085 112227 41113
rect 112261 41085 112289 41113
rect 112323 41085 112351 41113
rect 112137 41023 112165 41051
rect 112199 41023 112227 41051
rect 112261 41023 112289 41051
rect 112323 41023 112351 41051
rect 112137 40961 112165 40989
rect 112199 40961 112227 40989
rect 112261 40961 112289 40989
rect 112323 40961 112351 40989
rect 112137 32147 112165 32175
rect 112199 32147 112227 32175
rect 112261 32147 112289 32175
rect 112323 32147 112351 32175
rect 112137 32085 112165 32113
rect 112199 32085 112227 32113
rect 112261 32085 112289 32113
rect 112323 32085 112351 32113
rect 112137 32023 112165 32051
rect 112199 32023 112227 32051
rect 112261 32023 112289 32051
rect 112323 32023 112351 32051
rect 112137 31961 112165 31989
rect 112199 31961 112227 31989
rect 112261 31961 112289 31989
rect 112323 31961 112351 31989
rect 112137 23147 112165 23175
rect 112199 23147 112227 23175
rect 112261 23147 112289 23175
rect 112323 23147 112351 23175
rect 112137 23085 112165 23113
rect 112199 23085 112227 23113
rect 112261 23085 112289 23113
rect 112323 23085 112351 23113
rect 112137 23023 112165 23051
rect 112199 23023 112227 23051
rect 112261 23023 112289 23051
rect 112323 23023 112351 23051
rect 112137 22961 112165 22989
rect 112199 22961 112227 22989
rect 112261 22961 112289 22989
rect 112323 22961 112351 22989
rect 112137 14147 112165 14175
rect 112199 14147 112227 14175
rect 112261 14147 112289 14175
rect 112323 14147 112351 14175
rect 112137 14085 112165 14113
rect 112199 14085 112227 14113
rect 112261 14085 112289 14113
rect 112323 14085 112351 14113
rect 112137 14023 112165 14051
rect 112199 14023 112227 14051
rect 112261 14023 112289 14051
rect 112323 14023 112351 14051
rect 112137 13961 112165 13989
rect 112199 13961 112227 13989
rect 112261 13961 112289 13989
rect 112323 13961 112351 13989
rect 112137 5147 112165 5175
rect 112199 5147 112227 5175
rect 112261 5147 112289 5175
rect 112323 5147 112351 5175
rect 112137 5085 112165 5113
rect 112199 5085 112227 5113
rect 112261 5085 112289 5113
rect 112323 5085 112351 5113
rect 112137 5023 112165 5051
rect 112199 5023 112227 5051
rect 112261 5023 112289 5051
rect 112323 5023 112351 5051
rect 112137 4961 112165 4989
rect 112199 4961 112227 4989
rect 112261 4961 112289 4989
rect 112323 4961 112351 4989
rect 112137 -588 112165 -560
rect 112199 -588 112227 -560
rect 112261 -588 112289 -560
rect 112323 -588 112351 -560
rect 112137 -650 112165 -622
rect 112199 -650 112227 -622
rect 112261 -650 112289 -622
rect 112323 -650 112351 -622
rect 112137 -712 112165 -684
rect 112199 -712 112227 -684
rect 112261 -712 112289 -684
rect 112323 -712 112351 -684
rect 112137 -774 112165 -746
rect 112199 -774 112227 -746
rect 112261 -774 112289 -746
rect 112323 -774 112351 -746
rect 125637 92147 125665 92175
rect 125699 92147 125727 92175
rect 125761 92147 125789 92175
rect 125823 92147 125851 92175
rect 125637 92085 125665 92113
rect 125699 92085 125727 92113
rect 125761 92085 125789 92113
rect 125823 92085 125851 92113
rect 125637 92023 125665 92051
rect 125699 92023 125727 92051
rect 125761 92023 125789 92051
rect 125823 92023 125851 92051
rect 125637 91961 125665 91989
rect 125699 91961 125727 91989
rect 125761 91961 125789 91989
rect 125823 91961 125851 91989
rect 125637 83147 125665 83175
rect 125699 83147 125727 83175
rect 125761 83147 125789 83175
rect 125823 83147 125851 83175
rect 125637 83085 125665 83113
rect 125699 83085 125727 83113
rect 125761 83085 125789 83113
rect 125823 83085 125851 83113
rect 125637 83023 125665 83051
rect 125699 83023 125727 83051
rect 125761 83023 125789 83051
rect 125823 83023 125851 83051
rect 125637 82961 125665 82989
rect 125699 82961 125727 82989
rect 125761 82961 125789 82989
rect 125823 82961 125851 82989
rect 125637 74147 125665 74175
rect 125699 74147 125727 74175
rect 125761 74147 125789 74175
rect 125823 74147 125851 74175
rect 125637 74085 125665 74113
rect 125699 74085 125727 74113
rect 125761 74085 125789 74113
rect 125823 74085 125851 74113
rect 125637 74023 125665 74051
rect 125699 74023 125727 74051
rect 125761 74023 125789 74051
rect 125823 74023 125851 74051
rect 125637 73961 125665 73989
rect 125699 73961 125727 73989
rect 125761 73961 125789 73989
rect 125823 73961 125851 73989
rect 125637 65147 125665 65175
rect 125699 65147 125727 65175
rect 125761 65147 125789 65175
rect 125823 65147 125851 65175
rect 125637 65085 125665 65113
rect 125699 65085 125727 65113
rect 125761 65085 125789 65113
rect 125823 65085 125851 65113
rect 125637 65023 125665 65051
rect 125699 65023 125727 65051
rect 125761 65023 125789 65051
rect 125823 65023 125851 65051
rect 125637 64961 125665 64989
rect 125699 64961 125727 64989
rect 125761 64961 125789 64989
rect 125823 64961 125851 64989
rect 125637 56147 125665 56175
rect 125699 56147 125727 56175
rect 125761 56147 125789 56175
rect 125823 56147 125851 56175
rect 125637 56085 125665 56113
rect 125699 56085 125727 56113
rect 125761 56085 125789 56113
rect 125823 56085 125851 56113
rect 125637 56023 125665 56051
rect 125699 56023 125727 56051
rect 125761 56023 125789 56051
rect 125823 56023 125851 56051
rect 125637 55961 125665 55989
rect 125699 55961 125727 55989
rect 125761 55961 125789 55989
rect 125823 55961 125851 55989
rect 125637 47147 125665 47175
rect 125699 47147 125727 47175
rect 125761 47147 125789 47175
rect 125823 47147 125851 47175
rect 125637 47085 125665 47113
rect 125699 47085 125727 47113
rect 125761 47085 125789 47113
rect 125823 47085 125851 47113
rect 125637 47023 125665 47051
rect 125699 47023 125727 47051
rect 125761 47023 125789 47051
rect 125823 47023 125851 47051
rect 125637 46961 125665 46989
rect 125699 46961 125727 46989
rect 125761 46961 125789 46989
rect 125823 46961 125851 46989
rect 125637 38147 125665 38175
rect 125699 38147 125727 38175
rect 125761 38147 125789 38175
rect 125823 38147 125851 38175
rect 125637 38085 125665 38113
rect 125699 38085 125727 38113
rect 125761 38085 125789 38113
rect 125823 38085 125851 38113
rect 125637 38023 125665 38051
rect 125699 38023 125727 38051
rect 125761 38023 125789 38051
rect 125823 38023 125851 38051
rect 125637 37961 125665 37989
rect 125699 37961 125727 37989
rect 125761 37961 125789 37989
rect 125823 37961 125851 37989
rect 125637 29147 125665 29175
rect 125699 29147 125727 29175
rect 125761 29147 125789 29175
rect 125823 29147 125851 29175
rect 125637 29085 125665 29113
rect 125699 29085 125727 29113
rect 125761 29085 125789 29113
rect 125823 29085 125851 29113
rect 125637 29023 125665 29051
rect 125699 29023 125727 29051
rect 125761 29023 125789 29051
rect 125823 29023 125851 29051
rect 125637 28961 125665 28989
rect 125699 28961 125727 28989
rect 125761 28961 125789 28989
rect 125823 28961 125851 28989
rect 125637 20147 125665 20175
rect 125699 20147 125727 20175
rect 125761 20147 125789 20175
rect 125823 20147 125851 20175
rect 125637 20085 125665 20113
rect 125699 20085 125727 20113
rect 125761 20085 125789 20113
rect 125823 20085 125851 20113
rect 125637 20023 125665 20051
rect 125699 20023 125727 20051
rect 125761 20023 125789 20051
rect 125823 20023 125851 20051
rect 125637 19961 125665 19989
rect 125699 19961 125727 19989
rect 125761 19961 125789 19989
rect 125823 19961 125851 19989
rect 125637 11147 125665 11175
rect 125699 11147 125727 11175
rect 125761 11147 125789 11175
rect 125823 11147 125851 11175
rect 125637 11085 125665 11113
rect 125699 11085 125727 11113
rect 125761 11085 125789 11113
rect 125823 11085 125851 11113
rect 125637 11023 125665 11051
rect 125699 11023 125727 11051
rect 125761 11023 125789 11051
rect 125823 11023 125851 11051
rect 125637 10961 125665 10989
rect 125699 10961 125727 10989
rect 125761 10961 125789 10989
rect 125823 10961 125851 10989
rect 125637 2147 125665 2175
rect 125699 2147 125727 2175
rect 125761 2147 125789 2175
rect 125823 2147 125851 2175
rect 125637 2085 125665 2113
rect 125699 2085 125727 2113
rect 125761 2085 125789 2113
rect 125823 2085 125851 2113
rect 125637 2023 125665 2051
rect 125699 2023 125727 2051
rect 125761 2023 125789 2051
rect 125823 2023 125851 2051
rect 125637 1961 125665 1989
rect 125699 1961 125727 1989
rect 125761 1961 125789 1989
rect 125823 1961 125851 1989
rect 125637 -108 125665 -80
rect 125699 -108 125727 -80
rect 125761 -108 125789 -80
rect 125823 -108 125851 -80
rect 125637 -170 125665 -142
rect 125699 -170 125727 -142
rect 125761 -170 125789 -142
rect 125823 -170 125851 -142
rect 125637 -232 125665 -204
rect 125699 -232 125727 -204
rect 125761 -232 125789 -204
rect 125823 -232 125851 -204
rect 125637 -294 125665 -266
rect 125699 -294 125727 -266
rect 125761 -294 125789 -266
rect 125823 -294 125851 -266
rect 127497 95147 127525 95175
rect 127559 95147 127587 95175
rect 127621 95147 127649 95175
rect 127683 95147 127711 95175
rect 127497 95085 127525 95113
rect 127559 95085 127587 95113
rect 127621 95085 127649 95113
rect 127683 95085 127711 95113
rect 127497 95023 127525 95051
rect 127559 95023 127587 95051
rect 127621 95023 127649 95051
rect 127683 95023 127711 95051
rect 127497 94961 127525 94989
rect 127559 94961 127587 94989
rect 127621 94961 127649 94989
rect 127683 94961 127711 94989
rect 127497 86147 127525 86175
rect 127559 86147 127587 86175
rect 127621 86147 127649 86175
rect 127683 86147 127711 86175
rect 127497 86085 127525 86113
rect 127559 86085 127587 86113
rect 127621 86085 127649 86113
rect 127683 86085 127711 86113
rect 127497 86023 127525 86051
rect 127559 86023 127587 86051
rect 127621 86023 127649 86051
rect 127683 86023 127711 86051
rect 127497 85961 127525 85989
rect 127559 85961 127587 85989
rect 127621 85961 127649 85989
rect 127683 85961 127711 85989
rect 127497 77147 127525 77175
rect 127559 77147 127587 77175
rect 127621 77147 127649 77175
rect 127683 77147 127711 77175
rect 127497 77085 127525 77113
rect 127559 77085 127587 77113
rect 127621 77085 127649 77113
rect 127683 77085 127711 77113
rect 127497 77023 127525 77051
rect 127559 77023 127587 77051
rect 127621 77023 127649 77051
rect 127683 77023 127711 77051
rect 127497 76961 127525 76989
rect 127559 76961 127587 76989
rect 127621 76961 127649 76989
rect 127683 76961 127711 76989
rect 127497 68147 127525 68175
rect 127559 68147 127587 68175
rect 127621 68147 127649 68175
rect 127683 68147 127711 68175
rect 127497 68085 127525 68113
rect 127559 68085 127587 68113
rect 127621 68085 127649 68113
rect 127683 68085 127711 68113
rect 127497 68023 127525 68051
rect 127559 68023 127587 68051
rect 127621 68023 127649 68051
rect 127683 68023 127711 68051
rect 127497 67961 127525 67989
rect 127559 67961 127587 67989
rect 127621 67961 127649 67989
rect 127683 67961 127711 67989
rect 127497 59147 127525 59175
rect 127559 59147 127587 59175
rect 127621 59147 127649 59175
rect 127683 59147 127711 59175
rect 127497 59085 127525 59113
rect 127559 59085 127587 59113
rect 127621 59085 127649 59113
rect 127683 59085 127711 59113
rect 127497 59023 127525 59051
rect 127559 59023 127587 59051
rect 127621 59023 127649 59051
rect 127683 59023 127711 59051
rect 127497 58961 127525 58989
rect 127559 58961 127587 58989
rect 127621 58961 127649 58989
rect 127683 58961 127711 58989
rect 127497 50147 127525 50175
rect 127559 50147 127587 50175
rect 127621 50147 127649 50175
rect 127683 50147 127711 50175
rect 127497 50085 127525 50113
rect 127559 50085 127587 50113
rect 127621 50085 127649 50113
rect 127683 50085 127711 50113
rect 127497 50023 127525 50051
rect 127559 50023 127587 50051
rect 127621 50023 127649 50051
rect 127683 50023 127711 50051
rect 127497 49961 127525 49989
rect 127559 49961 127587 49989
rect 127621 49961 127649 49989
rect 127683 49961 127711 49989
rect 127497 41147 127525 41175
rect 127559 41147 127587 41175
rect 127621 41147 127649 41175
rect 127683 41147 127711 41175
rect 127497 41085 127525 41113
rect 127559 41085 127587 41113
rect 127621 41085 127649 41113
rect 127683 41085 127711 41113
rect 127497 41023 127525 41051
rect 127559 41023 127587 41051
rect 127621 41023 127649 41051
rect 127683 41023 127711 41051
rect 127497 40961 127525 40989
rect 127559 40961 127587 40989
rect 127621 40961 127649 40989
rect 127683 40961 127711 40989
rect 127497 32147 127525 32175
rect 127559 32147 127587 32175
rect 127621 32147 127649 32175
rect 127683 32147 127711 32175
rect 127497 32085 127525 32113
rect 127559 32085 127587 32113
rect 127621 32085 127649 32113
rect 127683 32085 127711 32113
rect 127497 32023 127525 32051
rect 127559 32023 127587 32051
rect 127621 32023 127649 32051
rect 127683 32023 127711 32051
rect 127497 31961 127525 31989
rect 127559 31961 127587 31989
rect 127621 31961 127649 31989
rect 127683 31961 127711 31989
rect 127497 23147 127525 23175
rect 127559 23147 127587 23175
rect 127621 23147 127649 23175
rect 127683 23147 127711 23175
rect 127497 23085 127525 23113
rect 127559 23085 127587 23113
rect 127621 23085 127649 23113
rect 127683 23085 127711 23113
rect 127497 23023 127525 23051
rect 127559 23023 127587 23051
rect 127621 23023 127649 23051
rect 127683 23023 127711 23051
rect 127497 22961 127525 22989
rect 127559 22961 127587 22989
rect 127621 22961 127649 22989
rect 127683 22961 127711 22989
rect 127497 14147 127525 14175
rect 127559 14147 127587 14175
rect 127621 14147 127649 14175
rect 127683 14147 127711 14175
rect 127497 14085 127525 14113
rect 127559 14085 127587 14113
rect 127621 14085 127649 14113
rect 127683 14085 127711 14113
rect 127497 14023 127525 14051
rect 127559 14023 127587 14051
rect 127621 14023 127649 14051
rect 127683 14023 127711 14051
rect 127497 13961 127525 13989
rect 127559 13961 127587 13989
rect 127621 13961 127649 13989
rect 127683 13961 127711 13989
rect 127497 5147 127525 5175
rect 127559 5147 127587 5175
rect 127621 5147 127649 5175
rect 127683 5147 127711 5175
rect 127497 5085 127525 5113
rect 127559 5085 127587 5113
rect 127621 5085 127649 5113
rect 127683 5085 127711 5113
rect 127497 5023 127525 5051
rect 127559 5023 127587 5051
rect 127621 5023 127649 5051
rect 127683 5023 127711 5051
rect 127497 4961 127525 4989
rect 127559 4961 127587 4989
rect 127621 4961 127649 4989
rect 127683 4961 127711 4989
rect 127497 -588 127525 -560
rect 127559 -588 127587 -560
rect 127621 -588 127649 -560
rect 127683 -588 127711 -560
rect 127497 -650 127525 -622
rect 127559 -650 127587 -622
rect 127621 -650 127649 -622
rect 127683 -650 127711 -622
rect 127497 -712 127525 -684
rect 127559 -712 127587 -684
rect 127621 -712 127649 -684
rect 127683 -712 127711 -684
rect 127497 -774 127525 -746
rect 127559 -774 127587 -746
rect 127621 -774 127649 -746
rect 127683 -774 127711 -746
rect 140997 92147 141025 92175
rect 141059 92147 141087 92175
rect 141121 92147 141149 92175
rect 141183 92147 141211 92175
rect 140997 92085 141025 92113
rect 141059 92085 141087 92113
rect 141121 92085 141149 92113
rect 141183 92085 141211 92113
rect 140997 92023 141025 92051
rect 141059 92023 141087 92051
rect 141121 92023 141149 92051
rect 141183 92023 141211 92051
rect 140997 91961 141025 91989
rect 141059 91961 141087 91989
rect 141121 91961 141149 91989
rect 141183 91961 141211 91989
rect 140997 83147 141025 83175
rect 141059 83147 141087 83175
rect 141121 83147 141149 83175
rect 141183 83147 141211 83175
rect 140997 83085 141025 83113
rect 141059 83085 141087 83113
rect 141121 83085 141149 83113
rect 141183 83085 141211 83113
rect 140997 83023 141025 83051
rect 141059 83023 141087 83051
rect 141121 83023 141149 83051
rect 141183 83023 141211 83051
rect 140997 82961 141025 82989
rect 141059 82961 141087 82989
rect 141121 82961 141149 82989
rect 141183 82961 141211 82989
rect 140997 74147 141025 74175
rect 141059 74147 141087 74175
rect 141121 74147 141149 74175
rect 141183 74147 141211 74175
rect 140997 74085 141025 74113
rect 141059 74085 141087 74113
rect 141121 74085 141149 74113
rect 141183 74085 141211 74113
rect 140997 74023 141025 74051
rect 141059 74023 141087 74051
rect 141121 74023 141149 74051
rect 141183 74023 141211 74051
rect 140997 73961 141025 73989
rect 141059 73961 141087 73989
rect 141121 73961 141149 73989
rect 141183 73961 141211 73989
rect 140997 65147 141025 65175
rect 141059 65147 141087 65175
rect 141121 65147 141149 65175
rect 141183 65147 141211 65175
rect 140997 65085 141025 65113
rect 141059 65085 141087 65113
rect 141121 65085 141149 65113
rect 141183 65085 141211 65113
rect 140997 65023 141025 65051
rect 141059 65023 141087 65051
rect 141121 65023 141149 65051
rect 141183 65023 141211 65051
rect 140997 64961 141025 64989
rect 141059 64961 141087 64989
rect 141121 64961 141149 64989
rect 141183 64961 141211 64989
rect 140997 56147 141025 56175
rect 141059 56147 141087 56175
rect 141121 56147 141149 56175
rect 141183 56147 141211 56175
rect 140997 56085 141025 56113
rect 141059 56085 141087 56113
rect 141121 56085 141149 56113
rect 141183 56085 141211 56113
rect 140997 56023 141025 56051
rect 141059 56023 141087 56051
rect 141121 56023 141149 56051
rect 141183 56023 141211 56051
rect 140997 55961 141025 55989
rect 141059 55961 141087 55989
rect 141121 55961 141149 55989
rect 141183 55961 141211 55989
rect 140997 47147 141025 47175
rect 141059 47147 141087 47175
rect 141121 47147 141149 47175
rect 141183 47147 141211 47175
rect 140997 47085 141025 47113
rect 141059 47085 141087 47113
rect 141121 47085 141149 47113
rect 141183 47085 141211 47113
rect 140997 47023 141025 47051
rect 141059 47023 141087 47051
rect 141121 47023 141149 47051
rect 141183 47023 141211 47051
rect 140997 46961 141025 46989
rect 141059 46961 141087 46989
rect 141121 46961 141149 46989
rect 141183 46961 141211 46989
rect 140997 38147 141025 38175
rect 141059 38147 141087 38175
rect 141121 38147 141149 38175
rect 141183 38147 141211 38175
rect 140997 38085 141025 38113
rect 141059 38085 141087 38113
rect 141121 38085 141149 38113
rect 141183 38085 141211 38113
rect 140997 38023 141025 38051
rect 141059 38023 141087 38051
rect 141121 38023 141149 38051
rect 141183 38023 141211 38051
rect 140997 37961 141025 37989
rect 141059 37961 141087 37989
rect 141121 37961 141149 37989
rect 141183 37961 141211 37989
rect 140997 29147 141025 29175
rect 141059 29147 141087 29175
rect 141121 29147 141149 29175
rect 141183 29147 141211 29175
rect 140997 29085 141025 29113
rect 141059 29085 141087 29113
rect 141121 29085 141149 29113
rect 141183 29085 141211 29113
rect 140997 29023 141025 29051
rect 141059 29023 141087 29051
rect 141121 29023 141149 29051
rect 141183 29023 141211 29051
rect 140997 28961 141025 28989
rect 141059 28961 141087 28989
rect 141121 28961 141149 28989
rect 141183 28961 141211 28989
rect 140997 20147 141025 20175
rect 141059 20147 141087 20175
rect 141121 20147 141149 20175
rect 141183 20147 141211 20175
rect 140997 20085 141025 20113
rect 141059 20085 141087 20113
rect 141121 20085 141149 20113
rect 141183 20085 141211 20113
rect 140997 20023 141025 20051
rect 141059 20023 141087 20051
rect 141121 20023 141149 20051
rect 141183 20023 141211 20051
rect 140997 19961 141025 19989
rect 141059 19961 141087 19989
rect 141121 19961 141149 19989
rect 141183 19961 141211 19989
rect 140997 11147 141025 11175
rect 141059 11147 141087 11175
rect 141121 11147 141149 11175
rect 141183 11147 141211 11175
rect 140997 11085 141025 11113
rect 141059 11085 141087 11113
rect 141121 11085 141149 11113
rect 141183 11085 141211 11113
rect 140997 11023 141025 11051
rect 141059 11023 141087 11051
rect 141121 11023 141149 11051
rect 141183 11023 141211 11051
rect 140997 10961 141025 10989
rect 141059 10961 141087 10989
rect 141121 10961 141149 10989
rect 141183 10961 141211 10989
rect 140997 2147 141025 2175
rect 141059 2147 141087 2175
rect 141121 2147 141149 2175
rect 141183 2147 141211 2175
rect 140997 2085 141025 2113
rect 141059 2085 141087 2113
rect 141121 2085 141149 2113
rect 141183 2085 141211 2113
rect 140997 2023 141025 2051
rect 141059 2023 141087 2051
rect 141121 2023 141149 2051
rect 141183 2023 141211 2051
rect 140997 1961 141025 1989
rect 141059 1961 141087 1989
rect 141121 1961 141149 1989
rect 141183 1961 141211 1989
rect 140997 -108 141025 -80
rect 141059 -108 141087 -80
rect 141121 -108 141149 -80
rect 141183 -108 141211 -80
rect 140997 -170 141025 -142
rect 141059 -170 141087 -142
rect 141121 -170 141149 -142
rect 141183 -170 141211 -142
rect 140997 -232 141025 -204
rect 141059 -232 141087 -204
rect 141121 -232 141149 -204
rect 141183 -232 141211 -204
rect 140997 -294 141025 -266
rect 141059 -294 141087 -266
rect 141121 -294 141149 -266
rect 141183 -294 141211 -266
rect 142857 95147 142885 95175
rect 142919 95147 142947 95175
rect 142981 95147 143009 95175
rect 143043 95147 143071 95175
rect 142857 95085 142885 95113
rect 142919 95085 142947 95113
rect 142981 95085 143009 95113
rect 143043 95085 143071 95113
rect 142857 95023 142885 95051
rect 142919 95023 142947 95051
rect 142981 95023 143009 95051
rect 143043 95023 143071 95051
rect 142857 94961 142885 94989
rect 142919 94961 142947 94989
rect 142981 94961 143009 94989
rect 143043 94961 143071 94989
rect 142857 86147 142885 86175
rect 142919 86147 142947 86175
rect 142981 86147 143009 86175
rect 143043 86147 143071 86175
rect 142857 86085 142885 86113
rect 142919 86085 142947 86113
rect 142981 86085 143009 86113
rect 143043 86085 143071 86113
rect 142857 86023 142885 86051
rect 142919 86023 142947 86051
rect 142981 86023 143009 86051
rect 143043 86023 143071 86051
rect 142857 85961 142885 85989
rect 142919 85961 142947 85989
rect 142981 85961 143009 85989
rect 143043 85961 143071 85989
rect 142857 77147 142885 77175
rect 142919 77147 142947 77175
rect 142981 77147 143009 77175
rect 143043 77147 143071 77175
rect 142857 77085 142885 77113
rect 142919 77085 142947 77113
rect 142981 77085 143009 77113
rect 143043 77085 143071 77113
rect 142857 77023 142885 77051
rect 142919 77023 142947 77051
rect 142981 77023 143009 77051
rect 143043 77023 143071 77051
rect 142857 76961 142885 76989
rect 142919 76961 142947 76989
rect 142981 76961 143009 76989
rect 143043 76961 143071 76989
rect 142857 68147 142885 68175
rect 142919 68147 142947 68175
rect 142981 68147 143009 68175
rect 143043 68147 143071 68175
rect 142857 68085 142885 68113
rect 142919 68085 142947 68113
rect 142981 68085 143009 68113
rect 143043 68085 143071 68113
rect 142857 68023 142885 68051
rect 142919 68023 142947 68051
rect 142981 68023 143009 68051
rect 143043 68023 143071 68051
rect 142857 67961 142885 67989
rect 142919 67961 142947 67989
rect 142981 67961 143009 67989
rect 143043 67961 143071 67989
rect 142857 59147 142885 59175
rect 142919 59147 142947 59175
rect 142981 59147 143009 59175
rect 143043 59147 143071 59175
rect 142857 59085 142885 59113
rect 142919 59085 142947 59113
rect 142981 59085 143009 59113
rect 143043 59085 143071 59113
rect 142857 59023 142885 59051
rect 142919 59023 142947 59051
rect 142981 59023 143009 59051
rect 143043 59023 143071 59051
rect 142857 58961 142885 58989
rect 142919 58961 142947 58989
rect 142981 58961 143009 58989
rect 143043 58961 143071 58989
rect 142857 50147 142885 50175
rect 142919 50147 142947 50175
rect 142981 50147 143009 50175
rect 143043 50147 143071 50175
rect 142857 50085 142885 50113
rect 142919 50085 142947 50113
rect 142981 50085 143009 50113
rect 143043 50085 143071 50113
rect 142857 50023 142885 50051
rect 142919 50023 142947 50051
rect 142981 50023 143009 50051
rect 143043 50023 143071 50051
rect 142857 49961 142885 49989
rect 142919 49961 142947 49989
rect 142981 49961 143009 49989
rect 143043 49961 143071 49989
rect 142857 41147 142885 41175
rect 142919 41147 142947 41175
rect 142981 41147 143009 41175
rect 143043 41147 143071 41175
rect 142857 41085 142885 41113
rect 142919 41085 142947 41113
rect 142981 41085 143009 41113
rect 143043 41085 143071 41113
rect 142857 41023 142885 41051
rect 142919 41023 142947 41051
rect 142981 41023 143009 41051
rect 143043 41023 143071 41051
rect 142857 40961 142885 40989
rect 142919 40961 142947 40989
rect 142981 40961 143009 40989
rect 143043 40961 143071 40989
rect 142857 32147 142885 32175
rect 142919 32147 142947 32175
rect 142981 32147 143009 32175
rect 143043 32147 143071 32175
rect 142857 32085 142885 32113
rect 142919 32085 142947 32113
rect 142981 32085 143009 32113
rect 143043 32085 143071 32113
rect 142857 32023 142885 32051
rect 142919 32023 142947 32051
rect 142981 32023 143009 32051
rect 143043 32023 143071 32051
rect 142857 31961 142885 31989
rect 142919 31961 142947 31989
rect 142981 31961 143009 31989
rect 143043 31961 143071 31989
rect 142857 23147 142885 23175
rect 142919 23147 142947 23175
rect 142981 23147 143009 23175
rect 143043 23147 143071 23175
rect 142857 23085 142885 23113
rect 142919 23085 142947 23113
rect 142981 23085 143009 23113
rect 143043 23085 143071 23113
rect 142857 23023 142885 23051
rect 142919 23023 142947 23051
rect 142981 23023 143009 23051
rect 143043 23023 143071 23051
rect 142857 22961 142885 22989
rect 142919 22961 142947 22989
rect 142981 22961 143009 22989
rect 143043 22961 143071 22989
rect 142857 14147 142885 14175
rect 142919 14147 142947 14175
rect 142981 14147 143009 14175
rect 143043 14147 143071 14175
rect 142857 14085 142885 14113
rect 142919 14085 142947 14113
rect 142981 14085 143009 14113
rect 143043 14085 143071 14113
rect 142857 14023 142885 14051
rect 142919 14023 142947 14051
rect 142981 14023 143009 14051
rect 143043 14023 143071 14051
rect 142857 13961 142885 13989
rect 142919 13961 142947 13989
rect 142981 13961 143009 13989
rect 143043 13961 143071 13989
rect 142857 5147 142885 5175
rect 142919 5147 142947 5175
rect 142981 5147 143009 5175
rect 143043 5147 143071 5175
rect 142857 5085 142885 5113
rect 142919 5085 142947 5113
rect 142981 5085 143009 5113
rect 143043 5085 143071 5113
rect 142857 5023 142885 5051
rect 142919 5023 142947 5051
rect 142981 5023 143009 5051
rect 143043 5023 143071 5051
rect 142857 4961 142885 4989
rect 142919 4961 142947 4989
rect 142981 4961 143009 4989
rect 143043 4961 143071 4989
rect 142857 -588 142885 -560
rect 142919 -588 142947 -560
rect 142981 -588 143009 -560
rect 143043 -588 143071 -560
rect 142857 -650 142885 -622
rect 142919 -650 142947 -622
rect 142981 -650 143009 -622
rect 143043 -650 143071 -622
rect 142857 -712 142885 -684
rect 142919 -712 142947 -684
rect 142981 -712 143009 -684
rect 143043 -712 143071 -684
rect 142857 -774 142885 -746
rect 142919 -774 142947 -746
rect 142981 -774 143009 -746
rect 143043 -774 143071 -746
rect 156357 92147 156385 92175
rect 156419 92147 156447 92175
rect 156481 92147 156509 92175
rect 156543 92147 156571 92175
rect 156357 92085 156385 92113
rect 156419 92085 156447 92113
rect 156481 92085 156509 92113
rect 156543 92085 156571 92113
rect 156357 92023 156385 92051
rect 156419 92023 156447 92051
rect 156481 92023 156509 92051
rect 156543 92023 156571 92051
rect 156357 91961 156385 91989
rect 156419 91961 156447 91989
rect 156481 91961 156509 91989
rect 156543 91961 156571 91989
rect 156357 83147 156385 83175
rect 156419 83147 156447 83175
rect 156481 83147 156509 83175
rect 156543 83147 156571 83175
rect 156357 83085 156385 83113
rect 156419 83085 156447 83113
rect 156481 83085 156509 83113
rect 156543 83085 156571 83113
rect 156357 83023 156385 83051
rect 156419 83023 156447 83051
rect 156481 83023 156509 83051
rect 156543 83023 156571 83051
rect 156357 82961 156385 82989
rect 156419 82961 156447 82989
rect 156481 82961 156509 82989
rect 156543 82961 156571 82989
rect 156357 74147 156385 74175
rect 156419 74147 156447 74175
rect 156481 74147 156509 74175
rect 156543 74147 156571 74175
rect 156357 74085 156385 74113
rect 156419 74085 156447 74113
rect 156481 74085 156509 74113
rect 156543 74085 156571 74113
rect 156357 74023 156385 74051
rect 156419 74023 156447 74051
rect 156481 74023 156509 74051
rect 156543 74023 156571 74051
rect 156357 73961 156385 73989
rect 156419 73961 156447 73989
rect 156481 73961 156509 73989
rect 156543 73961 156571 73989
rect 156357 65147 156385 65175
rect 156419 65147 156447 65175
rect 156481 65147 156509 65175
rect 156543 65147 156571 65175
rect 156357 65085 156385 65113
rect 156419 65085 156447 65113
rect 156481 65085 156509 65113
rect 156543 65085 156571 65113
rect 156357 65023 156385 65051
rect 156419 65023 156447 65051
rect 156481 65023 156509 65051
rect 156543 65023 156571 65051
rect 156357 64961 156385 64989
rect 156419 64961 156447 64989
rect 156481 64961 156509 64989
rect 156543 64961 156571 64989
rect 156357 56147 156385 56175
rect 156419 56147 156447 56175
rect 156481 56147 156509 56175
rect 156543 56147 156571 56175
rect 156357 56085 156385 56113
rect 156419 56085 156447 56113
rect 156481 56085 156509 56113
rect 156543 56085 156571 56113
rect 156357 56023 156385 56051
rect 156419 56023 156447 56051
rect 156481 56023 156509 56051
rect 156543 56023 156571 56051
rect 156357 55961 156385 55989
rect 156419 55961 156447 55989
rect 156481 55961 156509 55989
rect 156543 55961 156571 55989
rect 156357 47147 156385 47175
rect 156419 47147 156447 47175
rect 156481 47147 156509 47175
rect 156543 47147 156571 47175
rect 156357 47085 156385 47113
rect 156419 47085 156447 47113
rect 156481 47085 156509 47113
rect 156543 47085 156571 47113
rect 156357 47023 156385 47051
rect 156419 47023 156447 47051
rect 156481 47023 156509 47051
rect 156543 47023 156571 47051
rect 156357 46961 156385 46989
rect 156419 46961 156447 46989
rect 156481 46961 156509 46989
rect 156543 46961 156571 46989
rect 156357 38147 156385 38175
rect 156419 38147 156447 38175
rect 156481 38147 156509 38175
rect 156543 38147 156571 38175
rect 156357 38085 156385 38113
rect 156419 38085 156447 38113
rect 156481 38085 156509 38113
rect 156543 38085 156571 38113
rect 156357 38023 156385 38051
rect 156419 38023 156447 38051
rect 156481 38023 156509 38051
rect 156543 38023 156571 38051
rect 156357 37961 156385 37989
rect 156419 37961 156447 37989
rect 156481 37961 156509 37989
rect 156543 37961 156571 37989
rect 156357 29147 156385 29175
rect 156419 29147 156447 29175
rect 156481 29147 156509 29175
rect 156543 29147 156571 29175
rect 156357 29085 156385 29113
rect 156419 29085 156447 29113
rect 156481 29085 156509 29113
rect 156543 29085 156571 29113
rect 156357 29023 156385 29051
rect 156419 29023 156447 29051
rect 156481 29023 156509 29051
rect 156543 29023 156571 29051
rect 156357 28961 156385 28989
rect 156419 28961 156447 28989
rect 156481 28961 156509 28989
rect 156543 28961 156571 28989
rect 156357 20147 156385 20175
rect 156419 20147 156447 20175
rect 156481 20147 156509 20175
rect 156543 20147 156571 20175
rect 156357 20085 156385 20113
rect 156419 20085 156447 20113
rect 156481 20085 156509 20113
rect 156543 20085 156571 20113
rect 156357 20023 156385 20051
rect 156419 20023 156447 20051
rect 156481 20023 156509 20051
rect 156543 20023 156571 20051
rect 156357 19961 156385 19989
rect 156419 19961 156447 19989
rect 156481 19961 156509 19989
rect 156543 19961 156571 19989
rect 156357 11147 156385 11175
rect 156419 11147 156447 11175
rect 156481 11147 156509 11175
rect 156543 11147 156571 11175
rect 156357 11085 156385 11113
rect 156419 11085 156447 11113
rect 156481 11085 156509 11113
rect 156543 11085 156571 11113
rect 156357 11023 156385 11051
rect 156419 11023 156447 11051
rect 156481 11023 156509 11051
rect 156543 11023 156571 11051
rect 156357 10961 156385 10989
rect 156419 10961 156447 10989
rect 156481 10961 156509 10989
rect 156543 10961 156571 10989
rect 156357 2147 156385 2175
rect 156419 2147 156447 2175
rect 156481 2147 156509 2175
rect 156543 2147 156571 2175
rect 156357 2085 156385 2113
rect 156419 2085 156447 2113
rect 156481 2085 156509 2113
rect 156543 2085 156571 2113
rect 156357 2023 156385 2051
rect 156419 2023 156447 2051
rect 156481 2023 156509 2051
rect 156543 2023 156571 2051
rect 156357 1961 156385 1989
rect 156419 1961 156447 1989
rect 156481 1961 156509 1989
rect 156543 1961 156571 1989
rect 156357 -108 156385 -80
rect 156419 -108 156447 -80
rect 156481 -108 156509 -80
rect 156543 -108 156571 -80
rect 156357 -170 156385 -142
rect 156419 -170 156447 -142
rect 156481 -170 156509 -142
rect 156543 -170 156571 -142
rect 156357 -232 156385 -204
rect 156419 -232 156447 -204
rect 156481 -232 156509 -204
rect 156543 -232 156571 -204
rect 156357 -294 156385 -266
rect 156419 -294 156447 -266
rect 156481 -294 156509 -266
rect 156543 -294 156571 -266
rect 158217 95147 158245 95175
rect 158279 95147 158307 95175
rect 158341 95147 158369 95175
rect 158403 95147 158431 95175
rect 158217 95085 158245 95113
rect 158279 95085 158307 95113
rect 158341 95085 158369 95113
rect 158403 95085 158431 95113
rect 158217 95023 158245 95051
rect 158279 95023 158307 95051
rect 158341 95023 158369 95051
rect 158403 95023 158431 95051
rect 158217 94961 158245 94989
rect 158279 94961 158307 94989
rect 158341 94961 158369 94989
rect 158403 94961 158431 94989
rect 158217 86147 158245 86175
rect 158279 86147 158307 86175
rect 158341 86147 158369 86175
rect 158403 86147 158431 86175
rect 158217 86085 158245 86113
rect 158279 86085 158307 86113
rect 158341 86085 158369 86113
rect 158403 86085 158431 86113
rect 158217 86023 158245 86051
rect 158279 86023 158307 86051
rect 158341 86023 158369 86051
rect 158403 86023 158431 86051
rect 158217 85961 158245 85989
rect 158279 85961 158307 85989
rect 158341 85961 158369 85989
rect 158403 85961 158431 85989
rect 158217 77147 158245 77175
rect 158279 77147 158307 77175
rect 158341 77147 158369 77175
rect 158403 77147 158431 77175
rect 158217 77085 158245 77113
rect 158279 77085 158307 77113
rect 158341 77085 158369 77113
rect 158403 77085 158431 77113
rect 158217 77023 158245 77051
rect 158279 77023 158307 77051
rect 158341 77023 158369 77051
rect 158403 77023 158431 77051
rect 158217 76961 158245 76989
rect 158279 76961 158307 76989
rect 158341 76961 158369 76989
rect 158403 76961 158431 76989
rect 158217 68147 158245 68175
rect 158279 68147 158307 68175
rect 158341 68147 158369 68175
rect 158403 68147 158431 68175
rect 158217 68085 158245 68113
rect 158279 68085 158307 68113
rect 158341 68085 158369 68113
rect 158403 68085 158431 68113
rect 158217 68023 158245 68051
rect 158279 68023 158307 68051
rect 158341 68023 158369 68051
rect 158403 68023 158431 68051
rect 158217 67961 158245 67989
rect 158279 67961 158307 67989
rect 158341 67961 158369 67989
rect 158403 67961 158431 67989
rect 158217 59147 158245 59175
rect 158279 59147 158307 59175
rect 158341 59147 158369 59175
rect 158403 59147 158431 59175
rect 158217 59085 158245 59113
rect 158279 59085 158307 59113
rect 158341 59085 158369 59113
rect 158403 59085 158431 59113
rect 158217 59023 158245 59051
rect 158279 59023 158307 59051
rect 158341 59023 158369 59051
rect 158403 59023 158431 59051
rect 158217 58961 158245 58989
rect 158279 58961 158307 58989
rect 158341 58961 158369 58989
rect 158403 58961 158431 58989
rect 158217 50147 158245 50175
rect 158279 50147 158307 50175
rect 158341 50147 158369 50175
rect 158403 50147 158431 50175
rect 158217 50085 158245 50113
rect 158279 50085 158307 50113
rect 158341 50085 158369 50113
rect 158403 50085 158431 50113
rect 158217 50023 158245 50051
rect 158279 50023 158307 50051
rect 158341 50023 158369 50051
rect 158403 50023 158431 50051
rect 158217 49961 158245 49989
rect 158279 49961 158307 49989
rect 158341 49961 158369 49989
rect 158403 49961 158431 49989
rect 158217 41147 158245 41175
rect 158279 41147 158307 41175
rect 158341 41147 158369 41175
rect 158403 41147 158431 41175
rect 158217 41085 158245 41113
rect 158279 41085 158307 41113
rect 158341 41085 158369 41113
rect 158403 41085 158431 41113
rect 158217 41023 158245 41051
rect 158279 41023 158307 41051
rect 158341 41023 158369 41051
rect 158403 41023 158431 41051
rect 158217 40961 158245 40989
rect 158279 40961 158307 40989
rect 158341 40961 158369 40989
rect 158403 40961 158431 40989
rect 158217 32147 158245 32175
rect 158279 32147 158307 32175
rect 158341 32147 158369 32175
rect 158403 32147 158431 32175
rect 158217 32085 158245 32113
rect 158279 32085 158307 32113
rect 158341 32085 158369 32113
rect 158403 32085 158431 32113
rect 158217 32023 158245 32051
rect 158279 32023 158307 32051
rect 158341 32023 158369 32051
rect 158403 32023 158431 32051
rect 158217 31961 158245 31989
rect 158279 31961 158307 31989
rect 158341 31961 158369 31989
rect 158403 31961 158431 31989
rect 158217 23147 158245 23175
rect 158279 23147 158307 23175
rect 158341 23147 158369 23175
rect 158403 23147 158431 23175
rect 158217 23085 158245 23113
rect 158279 23085 158307 23113
rect 158341 23085 158369 23113
rect 158403 23085 158431 23113
rect 158217 23023 158245 23051
rect 158279 23023 158307 23051
rect 158341 23023 158369 23051
rect 158403 23023 158431 23051
rect 158217 22961 158245 22989
rect 158279 22961 158307 22989
rect 158341 22961 158369 22989
rect 158403 22961 158431 22989
rect 158217 14147 158245 14175
rect 158279 14147 158307 14175
rect 158341 14147 158369 14175
rect 158403 14147 158431 14175
rect 158217 14085 158245 14113
rect 158279 14085 158307 14113
rect 158341 14085 158369 14113
rect 158403 14085 158431 14113
rect 158217 14023 158245 14051
rect 158279 14023 158307 14051
rect 158341 14023 158369 14051
rect 158403 14023 158431 14051
rect 158217 13961 158245 13989
rect 158279 13961 158307 13989
rect 158341 13961 158369 13989
rect 158403 13961 158431 13989
rect 158217 5147 158245 5175
rect 158279 5147 158307 5175
rect 158341 5147 158369 5175
rect 158403 5147 158431 5175
rect 158217 5085 158245 5113
rect 158279 5085 158307 5113
rect 158341 5085 158369 5113
rect 158403 5085 158431 5113
rect 158217 5023 158245 5051
rect 158279 5023 158307 5051
rect 158341 5023 158369 5051
rect 158403 5023 158431 5051
rect 158217 4961 158245 4989
rect 158279 4961 158307 4989
rect 158341 4961 158369 4989
rect 158403 4961 158431 4989
rect 158217 -588 158245 -560
rect 158279 -588 158307 -560
rect 158341 -588 158369 -560
rect 158403 -588 158431 -560
rect 158217 -650 158245 -622
rect 158279 -650 158307 -622
rect 158341 -650 158369 -622
rect 158403 -650 158431 -622
rect 158217 -712 158245 -684
rect 158279 -712 158307 -684
rect 158341 -712 158369 -684
rect 158403 -712 158431 -684
rect 158217 -774 158245 -746
rect 158279 -774 158307 -746
rect 158341 -774 158369 -746
rect 158403 -774 158431 -746
rect 171717 92147 171745 92175
rect 171779 92147 171807 92175
rect 171841 92147 171869 92175
rect 171903 92147 171931 92175
rect 171717 92085 171745 92113
rect 171779 92085 171807 92113
rect 171841 92085 171869 92113
rect 171903 92085 171931 92113
rect 171717 92023 171745 92051
rect 171779 92023 171807 92051
rect 171841 92023 171869 92051
rect 171903 92023 171931 92051
rect 171717 91961 171745 91989
rect 171779 91961 171807 91989
rect 171841 91961 171869 91989
rect 171903 91961 171931 91989
rect 171717 83147 171745 83175
rect 171779 83147 171807 83175
rect 171841 83147 171869 83175
rect 171903 83147 171931 83175
rect 171717 83085 171745 83113
rect 171779 83085 171807 83113
rect 171841 83085 171869 83113
rect 171903 83085 171931 83113
rect 171717 83023 171745 83051
rect 171779 83023 171807 83051
rect 171841 83023 171869 83051
rect 171903 83023 171931 83051
rect 171717 82961 171745 82989
rect 171779 82961 171807 82989
rect 171841 82961 171869 82989
rect 171903 82961 171931 82989
rect 171717 74147 171745 74175
rect 171779 74147 171807 74175
rect 171841 74147 171869 74175
rect 171903 74147 171931 74175
rect 171717 74085 171745 74113
rect 171779 74085 171807 74113
rect 171841 74085 171869 74113
rect 171903 74085 171931 74113
rect 171717 74023 171745 74051
rect 171779 74023 171807 74051
rect 171841 74023 171869 74051
rect 171903 74023 171931 74051
rect 171717 73961 171745 73989
rect 171779 73961 171807 73989
rect 171841 73961 171869 73989
rect 171903 73961 171931 73989
rect 171717 65147 171745 65175
rect 171779 65147 171807 65175
rect 171841 65147 171869 65175
rect 171903 65147 171931 65175
rect 171717 65085 171745 65113
rect 171779 65085 171807 65113
rect 171841 65085 171869 65113
rect 171903 65085 171931 65113
rect 171717 65023 171745 65051
rect 171779 65023 171807 65051
rect 171841 65023 171869 65051
rect 171903 65023 171931 65051
rect 171717 64961 171745 64989
rect 171779 64961 171807 64989
rect 171841 64961 171869 64989
rect 171903 64961 171931 64989
rect 171717 56147 171745 56175
rect 171779 56147 171807 56175
rect 171841 56147 171869 56175
rect 171903 56147 171931 56175
rect 171717 56085 171745 56113
rect 171779 56085 171807 56113
rect 171841 56085 171869 56113
rect 171903 56085 171931 56113
rect 171717 56023 171745 56051
rect 171779 56023 171807 56051
rect 171841 56023 171869 56051
rect 171903 56023 171931 56051
rect 171717 55961 171745 55989
rect 171779 55961 171807 55989
rect 171841 55961 171869 55989
rect 171903 55961 171931 55989
rect 171717 47147 171745 47175
rect 171779 47147 171807 47175
rect 171841 47147 171869 47175
rect 171903 47147 171931 47175
rect 171717 47085 171745 47113
rect 171779 47085 171807 47113
rect 171841 47085 171869 47113
rect 171903 47085 171931 47113
rect 171717 47023 171745 47051
rect 171779 47023 171807 47051
rect 171841 47023 171869 47051
rect 171903 47023 171931 47051
rect 171717 46961 171745 46989
rect 171779 46961 171807 46989
rect 171841 46961 171869 46989
rect 171903 46961 171931 46989
rect 171717 38147 171745 38175
rect 171779 38147 171807 38175
rect 171841 38147 171869 38175
rect 171903 38147 171931 38175
rect 171717 38085 171745 38113
rect 171779 38085 171807 38113
rect 171841 38085 171869 38113
rect 171903 38085 171931 38113
rect 171717 38023 171745 38051
rect 171779 38023 171807 38051
rect 171841 38023 171869 38051
rect 171903 38023 171931 38051
rect 171717 37961 171745 37989
rect 171779 37961 171807 37989
rect 171841 37961 171869 37989
rect 171903 37961 171931 37989
rect 171717 29147 171745 29175
rect 171779 29147 171807 29175
rect 171841 29147 171869 29175
rect 171903 29147 171931 29175
rect 171717 29085 171745 29113
rect 171779 29085 171807 29113
rect 171841 29085 171869 29113
rect 171903 29085 171931 29113
rect 171717 29023 171745 29051
rect 171779 29023 171807 29051
rect 171841 29023 171869 29051
rect 171903 29023 171931 29051
rect 171717 28961 171745 28989
rect 171779 28961 171807 28989
rect 171841 28961 171869 28989
rect 171903 28961 171931 28989
rect 171717 20147 171745 20175
rect 171779 20147 171807 20175
rect 171841 20147 171869 20175
rect 171903 20147 171931 20175
rect 171717 20085 171745 20113
rect 171779 20085 171807 20113
rect 171841 20085 171869 20113
rect 171903 20085 171931 20113
rect 171717 20023 171745 20051
rect 171779 20023 171807 20051
rect 171841 20023 171869 20051
rect 171903 20023 171931 20051
rect 171717 19961 171745 19989
rect 171779 19961 171807 19989
rect 171841 19961 171869 19989
rect 171903 19961 171931 19989
rect 171717 11147 171745 11175
rect 171779 11147 171807 11175
rect 171841 11147 171869 11175
rect 171903 11147 171931 11175
rect 171717 11085 171745 11113
rect 171779 11085 171807 11113
rect 171841 11085 171869 11113
rect 171903 11085 171931 11113
rect 171717 11023 171745 11051
rect 171779 11023 171807 11051
rect 171841 11023 171869 11051
rect 171903 11023 171931 11051
rect 171717 10961 171745 10989
rect 171779 10961 171807 10989
rect 171841 10961 171869 10989
rect 171903 10961 171931 10989
rect 171717 2147 171745 2175
rect 171779 2147 171807 2175
rect 171841 2147 171869 2175
rect 171903 2147 171931 2175
rect 171717 2085 171745 2113
rect 171779 2085 171807 2113
rect 171841 2085 171869 2113
rect 171903 2085 171931 2113
rect 171717 2023 171745 2051
rect 171779 2023 171807 2051
rect 171841 2023 171869 2051
rect 171903 2023 171931 2051
rect 171717 1961 171745 1989
rect 171779 1961 171807 1989
rect 171841 1961 171869 1989
rect 171903 1961 171931 1989
rect 171717 -108 171745 -80
rect 171779 -108 171807 -80
rect 171841 -108 171869 -80
rect 171903 -108 171931 -80
rect 171717 -170 171745 -142
rect 171779 -170 171807 -142
rect 171841 -170 171869 -142
rect 171903 -170 171931 -142
rect 171717 -232 171745 -204
rect 171779 -232 171807 -204
rect 171841 -232 171869 -204
rect 171903 -232 171931 -204
rect 171717 -294 171745 -266
rect 171779 -294 171807 -266
rect 171841 -294 171869 -266
rect 171903 -294 171931 -266
rect 173577 95147 173605 95175
rect 173639 95147 173667 95175
rect 173701 95147 173729 95175
rect 173763 95147 173791 95175
rect 173577 95085 173605 95113
rect 173639 95085 173667 95113
rect 173701 95085 173729 95113
rect 173763 95085 173791 95113
rect 173577 95023 173605 95051
rect 173639 95023 173667 95051
rect 173701 95023 173729 95051
rect 173763 95023 173791 95051
rect 173577 94961 173605 94989
rect 173639 94961 173667 94989
rect 173701 94961 173729 94989
rect 173763 94961 173791 94989
rect 173577 86147 173605 86175
rect 173639 86147 173667 86175
rect 173701 86147 173729 86175
rect 173763 86147 173791 86175
rect 173577 86085 173605 86113
rect 173639 86085 173667 86113
rect 173701 86085 173729 86113
rect 173763 86085 173791 86113
rect 173577 86023 173605 86051
rect 173639 86023 173667 86051
rect 173701 86023 173729 86051
rect 173763 86023 173791 86051
rect 173577 85961 173605 85989
rect 173639 85961 173667 85989
rect 173701 85961 173729 85989
rect 173763 85961 173791 85989
rect 173577 77147 173605 77175
rect 173639 77147 173667 77175
rect 173701 77147 173729 77175
rect 173763 77147 173791 77175
rect 173577 77085 173605 77113
rect 173639 77085 173667 77113
rect 173701 77085 173729 77113
rect 173763 77085 173791 77113
rect 173577 77023 173605 77051
rect 173639 77023 173667 77051
rect 173701 77023 173729 77051
rect 173763 77023 173791 77051
rect 173577 76961 173605 76989
rect 173639 76961 173667 76989
rect 173701 76961 173729 76989
rect 173763 76961 173791 76989
rect 173577 68147 173605 68175
rect 173639 68147 173667 68175
rect 173701 68147 173729 68175
rect 173763 68147 173791 68175
rect 173577 68085 173605 68113
rect 173639 68085 173667 68113
rect 173701 68085 173729 68113
rect 173763 68085 173791 68113
rect 173577 68023 173605 68051
rect 173639 68023 173667 68051
rect 173701 68023 173729 68051
rect 173763 68023 173791 68051
rect 173577 67961 173605 67989
rect 173639 67961 173667 67989
rect 173701 67961 173729 67989
rect 173763 67961 173791 67989
rect 173577 59147 173605 59175
rect 173639 59147 173667 59175
rect 173701 59147 173729 59175
rect 173763 59147 173791 59175
rect 173577 59085 173605 59113
rect 173639 59085 173667 59113
rect 173701 59085 173729 59113
rect 173763 59085 173791 59113
rect 173577 59023 173605 59051
rect 173639 59023 173667 59051
rect 173701 59023 173729 59051
rect 173763 59023 173791 59051
rect 173577 58961 173605 58989
rect 173639 58961 173667 58989
rect 173701 58961 173729 58989
rect 173763 58961 173791 58989
rect 173577 50147 173605 50175
rect 173639 50147 173667 50175
rect 173701 50147 173729 50175
rect 173763 50147 173791 50175
rect 173577 50085 173605 50113
rect 173639 50085 173667 50113
rect 173701 50085 173729 50113
rect 173763 50085 173791 50113
rect 173577 50023 173605 50051
rect 173639 50023 173667 50051
rect 173701 50023 173729 50051
rect 173763 50023 173791 50051
rect 173577 49961 173605 49989
rect 173639 49961 173667 49989
rect 173701 49961 173729 49989
rect 173763 49961 173791 49989
rect 173577 41147 173605 41175
rect 173639 41147 173667 41175
rect 173701 41147 173729 41175
rect 173763 41147 173791 41175
rect 173577 41085 173605 41113
rect 173639 41085 173667 41113
rect 173701 41085 173729 41113
rect 173763 41085 173791 41113
rect 173577 41023 173605 41051
rect 173639 41023 173667 41051
rect 173701 41023 173729 41051
rect 173763 41023 173791 41051
rect 173577 40961 173605 40989
rect 173639 40961 173667 40989
rect 173701 40961 173729 40989
rect 173763 40961 173791 40989
rect 173577 32147 173605 32175
rect 173639 32147 173667 32175
rect 173701 32147 173729 32175
rect 173763 32147 173791 32175
rect 173577 32085 173605 32113
rect 173639 32085 173667 32113
rect 173701 32085 173729 32113
rect 173763 32085 173791 32113
rect 173577 32023 173605 32051
rect 173639 32023 173667 32051
rect 173701 32023 173729 32051
rect 173763 32023 173791 32051
rect 173577 31961 173605 31989
rect 173639 31961 173667 31989
rect 173701 31961 173729 31989
rect 173763 31961 173791 31989
rect 173577 23147 173605 23175
rect 173639 23147 173667 23175
rect 173701 23147 173729 23175
rect 173763 23147 173791 23175
rect 173577 23085 173605 23113
rect 173639 23085 173667 23113
rect 173701 23085 173729 23113
rect 173763 23085 173791 23113
rect 173577 23023 173605 23051
rect 173639 23023 173667 23051
rect 173701 23023 173729 23051
rect 173763 23023 173791 23051
rect 173577 22961 173605 22989
rect 173639 22961 173667 22989
rect 173701 22961 173729 22989
rect 173763 22961 173791 22989
rect 173577 14147 173605 14175
rect 173639 14147 173667 14175
rect 173701 14147 173729 14175
rect 173763 14147 173791 14175
rect 173577 14085 173605 14113
rect 173639 14085 173667 14113
rect 173701 14085 173729 14113
rect 173763 14085 173791 14113
rect 173577 14023 173605 14051
rect 173639 14023 173667 14051
rect 173701 14023 173729 14051
rect 173763 14023 173791 14051
rect 173577 13961 173605 13989
rect 173639 13961 173667 13989
rect 173701 13961 173729 13989
rect 173763 13961 173791 13989
rect 173577 5147 173605 5175
rect 173639 5147 173667 5175
rect 173701 5147 173729 5175
rect 173763 5147 173791 5175
rect 173577 5085 173605 5113
rect 173639 5085 173667 5113
rect 173701 5085 173729 5113
rect 173763 5085 173791 5113
rect 173577 5023 173605 5051
rect 173639 5023 173667 5051
rect 173701 5023 173729 5051
rect 173763 5023 173791 5051
rect 173577 4961 173605 4989
rect 173639 4961 173667 4989
rect 173701 4961 173729 4989
rect 173763 4961 173791 4989
rect 173577 -588 173605 -560
rect 173639 -588 173667 -560
rect 173701 -588 173729 -560
rect 173763 -588 173791 -560
rect 173577 -650 173605 -622
rect 173639 -650 173667 -622
rect 173701 -650 173729 -622
rect 173763 -650 173791 -622
rect 173577 -712 173605 -684
rect 173639 -712 173667 -684
rect 173701 -712 173729 -684
rect 173763 -712 173791 -684
rect 173577 -774 173605 -746
rect 173639 -774 173667 -746
rect 173701 -774 173729 -746
rect 173763 -774 173791 -746
rect 187077 92147 187105 92175
rect 187139 92147 187167 92175
rect 187201 92147 187229 92175
rect 187263 92147 187291 92175
rect 187077 92085 187105 92113
rect 187139 92085 187167 92113
rect 187201 92085 187229 92113
rect 187263 92085 187291 92113
rect 187077 92023 187105 92051
rect 187139 92023 187167 92051
rect 187201 92023 187229 92051
rect 187263 92023 187291 92051
rect 187077 91961 187105 91989
rect 187139 91961 187167 91989
rect 187201 91961 187229 91989
rect 187263 91961 187291 91989
rect 187077 83147 187105 83175
rect 187139 83147 187167 83175
rect 187201 83147 187229 83175
rect 187263 83147 187291 83175
rect 187077 83085 187105 83113
rect 187139 83085 187167 83113
rect 187201 83085 187229 83113
rect 187263 83085 187291 83113
rect 187077 83023 187105 83051
rect 187139 83023 187167 83051
rect 187201 83023 187229 83051
rect 187263 83023 187291 83051
rect 187077 82961 187105 82989
rect 187139 82961 187167 82989
rect 187201 82961 187229 82989
rect 187263 82961 187291 82989
rect 187077 74147 187105 74175
rect 187139 74147 187167 74175
rect 187201 74147 187229 74175
rect 187263 74147 187291 74175
rect 187077 74085 187105 74113
rect 187139 74085 187167 74113
rect 187201 74085 187229 74113
rect 187263 74085 187291 74113
rect 187077 74023 187105 74051
rect 187139 74023 187167 74051
rect 187201 74023 187229 74051
rect 187263 74023 187291 74051
rect 187077 73961 187105 73989
rect 187139 73961 187167 73989
rect 187201 73961 187229 73989
rect 187263 73961 187291 73989
rect 187077 65147 187105 65175
rect 187139 65147 187167 65175
rect 187201 65147 187229 65175
rect 187263 65147 187291 65175
rect 187077 65085 187105 65113
rect 187139 65085 187167 65113
rect 187201 65085 187229 65113
rect 187263 65085 187291 65113
rect 187077 65023 187105 65051
rect 187139 65023 187167 65051
rect 187201 65023 187229 65051
rect 187263 65023 187291 65051
rect 187077 64961 187105 64989
rect 187139 64961 187167 64989
rect 187201 64961 187229 64989
rect 187263 64961 187291 64989
rect 187077 56147 187105 56175
rect 187139 56147 187167 56175
rect 187201 56147 187229 56175
rect 187263 56147 187291 56175
rect 187077 56085 187105 56113
rect 187139 56085 187167 56113
rect 187201 56085 187229 56113
rect 187263 56085 187291 56113
rect 187077 56023 187105 56051
rect 187139 56023 187167 56051
rect 187201 56023 187229 56051
rect 187263 56023 187291 56051
rect 187077 55961 187105 55989
rect 187139 55961 187167 55989
rect 187201 55961 187229 55989
rect 187263 55961 187291 55989
rect 187077 47147 187105 47175
rect 187139 47147 187167 47175
rect 187201 47147 187229 47175
rect 187263 47147 187291 47175
rect 187077 47085 187105 47113
rect 187139 47085 187167 47113
rect 187201 47085 187229 47113
rect 187263 47085 187291 47113
rect 187077 47023 187105 47051
rect 187139 47023 187167 47051
rect 187201 47023 187229 47051
rect 187263 47023 187291 47051
rect 187077 46961 187105 46989
rect 187139 46961 187167 46989
rect 187201 46961 187229 46989
rect 187263 46961 187291 46989
rect 187077 38147 187105 38175
rect 187139 38147 187167 38175
rect 187201 38147 187229 38175
rect 187263 38147 187291 38175
rect 187077 38085 187105 38113
rect 187139 38085 187167 38113
rect 187201 38085 187229 38113
rect 187263 38085 187291 38113
rect 187077 38023 187105 38051
rect 187139 38023 187167 38051
rect 187201 38023 187229 38051
rect 187263 38023 187291 38051
rect 187077 37961 187105 37989
rect 187139 37961 187167 37989
rect 187201 37961 187229 37989
rect 187263 37961 187291 37989
rect 187077 29147 187105 29175
rect 187139 29147 187167 29175
rect 187201 29147 187229 29175
rect 187263 29147 187291 29175
rect 187077 29085 187105 29113
rect 187139 29085 187167 29113
rect 187201 29085 187229 29113
rect 187263 29085 187291 29113
rect 187077 29023 187105 29051
rect 187139 29023 187167 29051
rect 187201 29023 187229 29051
rect 187263 29023 187291 29051
rect 187077 28961 187105 28989
rect 187139 28961 187167 28989
rect 187201 28961 187229 28989
rect 187263 28961 187291 28989
rect 187077 20147 187105 20175
rect 187139 20147 187167 20175
rect 187201 20147 187229 20175
rect 187263 20147 187291 20175
rect 187077 20085 187105 20113
rect 187139 20085 187167 20113
rect 187201 20085 187229 20113
rect 187263 20085 187291 20113
rect 187077 20023 187105 20051
rect 187139 20023 187167 20051
rect 187201 20023 187229 20051
rect 187263 20023 187291 20051
rect 187077 19961 187105 19989
rect 187139 19961 187167 19989
rect 187201 19961 187229 19989
rect 187263 19961 187291 19989
rect 187077 11147 187105 11175
rect 187139 11147 187167 11175
rect 187201 11147 187229 11175
rect 187263 11147 187291 11175
rect 187077 11085 187105 11113
rect 187139 11085 187167 11113
rect 187201 11085 187229 11113
rect 187263 11085 187291 11113
rect 187077 11023 187105 11051
rect 187139 11023 187167 11051
rect 187201 11023 187229 11051
rect 187263 11023 187291 11051
rect 187077 10961 187105 10989
rect 187139 10961 187167 10989
rect 187201 10961 187229 10989
rect 187263 10961 187291 10989
rect 187077 2147 187105 2175
rect 187139 2147 187167 2175
rect 187201 2147 187229 2175
rect 187263 2147 187291 2175
rect 187077 2085 187105 2113
rect 187139 2085 187167 2113
rect 187201 2085 187229 2113
rect 187263 2085 187291 2113
rect 187077 2023 187105 2051
rect 187139 2023 187167 2051
rect 187201 2023 187229 2051
rect 187263 2023 187291 2051
rect 187077 1961 187105 1989
rect 187139 1961 187167 1989
rect 187201 1961 187229 1989
rect 187263 1961 187291 1989
rect 187077 -108 187105 -80
rect 187139 -108 187167 -80
rect 187201 -108 187229 -80
rect 187263 -108 187291 -80
rect 187077 -170 187105 -142
rect 187139 -170 187167 -142
rect 187201 -170 187229 -142
rect 187263 -170 187291 -142
rect 187077 -232 187105 -204
rect 187139 -232 187167 -204
rect 187201 -232 187229 -204
rect 187263 -232 187291 -204
rect 187077 -294 187105 -266
rect 187139 -294 187167 -266
rect 187201 -294 187229 -266
rect 187263 -294 187291 -266
rect 188937 95147 188965 95175
rect 188999 95147 189027 95175
rect 189061 95147 189089 95175
rect 189123 95147 189151 95175
rect 188937 95085 188965 95113
rect 188999 95085 189027 95113
rect 189061 95085 189089 95113
rect 189123 95085 189151 95113
rect 188937 95023 188965 95051
rect 188999 95023 189027 95051
rect 189061 95023 189089 95051
rect 189123 95023 189151 95051
rect 188937 94961 188965 94989
rect 188999 94961 189027 94989
rect 189061 94961 189089 94989
rect 189123 94961 189151 94989
rect 188937 86147 188965 86175
rect 188999 86147 189027 86175
rect 189061 86147 189089 86175
rect 189123 86147 189151 86175
rect 188937 86085 188965 86113
rect 188999 86085 189027 86113
rect 189061 86085 189089 86113
rect 189123 86085 189151 86113
rect 188937 86023 188965 86051
rect 188999 86023 189027 86051
rect 189061 86023 189089 86051
rect 189123 86023 189151 86051
rect 188937 85961 188965 85989
rect 188999 85961 189027 85989
rect 189061 85961 189089 85989
rect 189123 85961 189151 85989
rect 188937 77147 188965 77175
rect 188999 77147 189027 77175
rect 189061 77147 189089 77175
rect 189123 77147 189151 77175
rect 188937 77085 188965 77113
rect 188999 77085 189027 77113
rect 189061 77085 189089 77113
rect 189123 77085 189151 77113
rect 188937 77023 188965 77051
rect 188999 77023 189027 77051
rect 189061 77023 189089 77051
rect 189123 77023 189151 77051
rect 188937 76961 188965 76989
rect 188999 76961 189027 76989
rect 189061 76961 189089 76989
rect 189123 76961 189151 76989
rect 188937 68147 188965 68175
rect 188999 68147 189027 68175
rect 189061 68147 189089 68175
rect 189123 68147 189151 68175
rect 188937 68085 188965 68113
rect 188999 68085 189027 68113
rect 189061 68085 189089 68113
rect 189123 68085 189151 68113
rect 188937 68023 188965 68051
rect 188999 68023 189027 68051
rect 189061 68023 189089 68051
rect 189123 68023 189151 68051
rect 188937 67961 188965 67989
rect 188999 67961 189027 67989
rect 189061 67961 189089 67989
rect 189123 67961 189151 67989
rect 188937 59147 188965 59175
rect 188999 59147 189027 59175
rect 189061 59147 189089 59175
rect 189123 59147 189151 59175
rect 188937 59085 188965 59113
rect 188999 59085 189027 59113
rect 189061 59085 189089 59113
rect 189123 59085 189151 59113
rect 188937 59023 188965 59051
rect 188999 59023 189027 59051
rect 189061 59023 189089 59051
rect 189123 59023 189151 59051
rect 188937 58961 188965 58989
rect 188999 58961 189027 58989
rect 189061 58961 189089 58989
rect 189123 58961 189151 58989
rect 188937 50147 188965 50175
rect 188999 50147 189027 50175
rect 189061 50147 189089 50175
rect 189123 50147 189151 50175
rect 188937 50085 188965 50113
rect 188999 50085 189027 50113
rect 189061 50085 189089 50113
rect 189123 50085 189151 50113
rect 188937 50023 188965 50051
rect 188999 50023 189027 50051
rect 189061 50023 189089 50051
rect 189123 50023 189151 50051
rect 188937 49961 188965 49989
rect 188999 49961 189027 49989
rect 189061 49961 189089 49989
rect 189123 49961 189151 49989
rect 188937 41147 188965 41175
rect 188999 41147 189027 41175
rect 189061 41147 189089 41175
rect 189123 41147 189151 41175
rect 188937 41085 188965 41113
rect 188999 41085 189027 41113
rect 189061 41085 189089 41113
rect 189123 41085 189151 41113
rect 188937 41023 188965 41051
rect 188999 41023 189027 41051
rect 189061 41023 189089 41051
rect 189123 41023 189151 41051
rect 188937 40961 188965 40989
rect 188999 40961 189027 40989
rect 189061 40961 189089 40989
rect 189123 40961 189151 40989
rect 188937 32147 188965 32175
rect 188999 32147 189027 32175
rect 189061 32147 189089 32175
rect 189123 32147 189151 32175
rect 188937 32085 188965 32113
rect 188999 32085 189027 32113
rect 189061 32085 189089 32113
rect 189123 32085 189151 32113
rect 188937 32023 188965 32051
rect 188999 32023 189027 32051
rect 189061 32023 189089 32051
rect 189123 32023 189151 32051
rect 188937 31961 188965 31989
rect 188999 31961 189027 31989
rect 189061 31961 189089 31989
rect 189123 31961 189151 31989
rect 188937 23147 188965 23175
rect 188999 23147 189027 23175
rect 189061 23147 189089 23175
rect 189123 23147 189151 23175
rect 188937 23085 188965 23113
rect 188999 23085 189027 23113
rect 189061 23085 189089 23113
rect 189123 23085 189151 23113
rect 188937 23023 188965 23051
rect 188999 23023 189027 23051
rect 189061 23023 189089 23051
rect 189123 23023 189151 23051
rect 188937 22961 188965 22989
rect 188999 22961 189027 22989
rect 189061 22961 189089 22989
rect 189123 22961 189151 22989
rect 188937 14147 188965 14175
rect 188999 14147 189027 14175
rect 189061 14147 189089 14175
rect 189123 14147 189151 14175
rect 188937 14085 188965 14113
rect 188999 14085 189027 14113
rect 189061 14085 189089 14113
rect 189123 14085 189151 14113
rect 188937 14023 188965 14051
rect 188999 14023 189027 14051
rect 189061 14023 189089 14051
rect 189123 14023 189151 14051
rect 188937 13961 188965 13989
rect 188999 13961 189027 13989
rect 189061 13961 189089 13989
rect 189123 13961 189151 13989
rect 188937 5147 188965 5175
rect 188999 5147 189027 5175
rect 189061 5147 189089 5175
rect 189123 5147 189151 5175
rect 188937 5085 188965 5113
rect 188999 5085 189027 5113
rect 189061 5085 189089 5113
rect 189123 5085 189151 5113
rect 188937 5023 188965 5051
rect 188999 5023 189027 5051
rect 189061 5023 189089 5051
rect 189123 5023 189151 5051
rect 188937 4961 188965 4989
rect 188999 4961 189027 4989
rect 189061 4961 189089 4989
rect 189123 4961 189151 4989
rect 188937 -588 188965 -560
rect 188999 -588 189027 -560
rect 189061 -588 189089 -560
rect 189123 -588 189151 -560
rect 188937 -650 188965 -622
rect 188999 -650 189027 -622
rect 189061 -650 189089 -622
rect 189123 -650 189151 -622
rect 188937 -712 188965 -684
rect 188999 -712 189027 -684
rect 189061 -712 189089 -684
rect 189123 -712 189151 -684
rect 188937 -774 188965 -746
rect 188999 -774 189027 -746
rect 189061 -774 189089 -746
rect 189123 -774 189151 -746
rect 202437 92147 202465 92175
rect 202499 92147 202527 92175
rect 202561 92147 202589 92175
rect 202623 92147 202651 92175
rect 202437 92085 202465 92113
rect 202499 92085 202527 92113
rect 202561 92085 202589 92113
rect 202623 92085 202651 92113
rect 202437 92023 202465 92051
rect 202499 92023 202527 92051
rect 202561 92023 202589 92051
rect 202623 92023 202651 92051
rect 202437 91961 202465 91989
rect 202499 91961 202527 91989
rect 202561 91961 202589 91989
rect 202623 91961 202651 91989
rect 202437 83147 202465 83175
rect 202499 83147 202527 83175
rect 202561 83147 202589 83175
rect 202623 83147 202651 83175
rect 202437 83085 202465 83113
rect 202499 83085 202527 83113
rect 202561 83085 202589 83113
rect 202623 83085 202651 83113
rect 202437 83023 202465 83051
rect 202499 83023 202527 83051
rect 202561 83023 202589 83051
rect 202623 83023 202651 83051
rect 202437 82961 202465 82989
rect 202499 82961 202527 82989
rect 202561 82961 202589 82989
rect 202623 82961 202651 82989
rect 202437 74147 202465 74175
rect 202499 74147 202527 74175
rect 202561 74147 202589 74175
rect 202623 74147 202651 74175
rect 202437 74085 202465 74113
rect 202499 74085 202527 74113
rect 202561 74085 202589 74113
rect 202623 74085 202651 74113
rect 202437 74023 202465 74051
rect 202499 74023 202527 74051
rect 202561 74023 202589 74051
rect 202623 74023 202651 74051
rect 202437 73961 202465 73989
rect 202499 73961 202527 73989
rect 202561 73961 202589 73989
rect 202623 73961 202651 73989
rect 202437 65147 202465 65175
rect 202499 65147 202527 65175
rect 202561 65147 202589 65175
rect 202623 65147 202651 65175
rect 202437 65085 202465 65113
rect 202499 65085 202527 65113
rect 202561 65085 202589 65113
rect 202623 65085 202651 65113
rect 202437 65023 202465 65051
rect 202499 65023 202527 65051
rect 202561 65023 202589 65051
rect 202623 65023 202651 65051
rect 202437 64961 202465 64989
rect 202499 64961 202527 64989
rect 202561 64961 202589 64989
rect 202623 64961 202651 64989
rect 202437 56147 202465 56175
rect 202499 56147 202527 56175
rect 202561 56147 202589 56175
rect 202623 56147 202651 56175
rect 202437 56085 202465 56113
rect 202499 56085 202527 56113
rect 202561 56085 202589 56113
rect 202623 56085 202651 56113
rect 202437 56023 202465 56051
rect 202499 56023 202527 56051
rect 202561 56023 202589 56051
rect 202623 56023 202651 56051
rect 202437 55961 202465 55989
rect 202499 55961 202527 55989
rect 202561 55961 202589 55989
rect 202623 55961 202651 55989
rect 202437 47147 202465 47175
rect 202499 47147 202527 47175
rect 202561 47147 202589 47175
rect 202623 47147 202651 47175
rect 202437 47085 202465 47113
rect 202499 47085 202527 47113
rect 202561 47085 202589 47113
rect 202623 47085 202651 47113
rect 202437 47023 202465 47051
rect 202499 47023 202527 47051
rect 202561 47023 202589 47051
rect 202623 47023 202651 47051
rect 202437 46961 202465 46989
rect 202499 46961 202527 46989
rect 202561 46961 202589 46989
rect 202623 46961 202651 46989
rect 202437 38147 202465 38175
rect 202499 38147 202527 38175
rect 202561 38147 202589 38175
rect 202623 38147 202651 38175
rect 202437 38085 202465 38113
rect 202499 38085 202527 38113
rect 202561 38085 202589 38113
rect 202623 38085 202651 38113
rect 202437 38023 202465 38051
rect 202499 38023 202527 38051
rect 202561 38023 202589 38051
rect 202623 38023 202651 38051
rect 202437 37961 202465 37989
rect 202499 37961 202527 37989
rect 202561 37961 202589 37989
rect 202623 37961 202651 37989
rect 202437 29147 202465 29175
rect 202499 29147 202527 29175
rect 202561 29147 202589 29175
rect 202623 29147 202651 29175
rect 202437 29085 202465 29113
rect 202499 29085 202527 29113
rect 202561 29085 202589 29113
rect 202623 29085 202651 29113
rect 202437 29023 202465 29051
rect 202499 29023 202527 29051
rect 202561 29023 202589 29051
rect 202623 29023 202651 29051
rect 202437 28961 202465 28989
rect 202499 28961 202527 28989
rect 202561 28961 202589 28989
rect 202623 28961 202651 28989
rect 202437 20147 202465 20175
rect 202499 20147 202527 20175
rect 202561 20147 202589 20175
rect 202623 20147 202651 20175
rect 202437 20085 202465 20113
rect 202499 20085 202527 20113
rect 202561 20085 202589 20113
rect 202623 20085 202651 20113
rect 202437 20023 202465 20051
rect 202499 20023 202527 20051
rect 202561 20023 202589 20051
rect 202623 20023 202651 20051
rect 202437 19961 202465 19989
rect 202499 19961 202527 19989
rect 202561 19961 202589 19989
rect 202623 19961 202651 19989
rect 202437 11147 202465 11175
rect 202499 11147 202527 11175
rect 202561 11147 202589 11175
rect 202623 11147 202651 11175
rect 202437 11085 202465 11113
rect 202499 11085 202527 11113
rect 202561 11085 202589 11113
rect 202623 11085 202651 11113
rect 202437 11023 202465 11051
rect 202499 11023 202527 11051
rect 202561 11023 202589 11051
rect 202623 11023 202651 11051
rect 202437 10961 202465 10989
rect 202499 10961 202527 10989
rect 202561 10961 202589 10989
rect 202623 10961 202651 10989
rect 202437 2147 202465 2175
rect 202499 2147 202527 2175
rect 202561 2147 202589 2175
rect 202623 2147 202651 2175
rect 202437 2085 202465 2113
rect 202499 2085 202527 2113
rect 202561 2085 202589 2113
rect 202623 2085 202651 2113
rect 202437 2023 202465 2051
rect 202499 2023 202527 2051
rect 202561 2023 202589 2051
rect 202623 2023 202651 2051
rect 202437 1961 202465 1989
rect 202499 1961 202527 1989
rect 202561 1961 202589 1989
rect 202623 1961 202651 1989
rect 202437 -108 202465 -80
rect 202499 -108 202527 -80
rect 202561 -108 202589 -80
rect 202623 -108 202651 -80
rect 202437 -170 202465 -142
rect 202499 -170 202527 -142
rect 202561 -170 202589 -142
rect 202623 -170 202651 -142
rect 202437 -232 202465 -204
rect 202499 -232 202527 -204
rect 202561 -232 202589 -204
rect 202623 -232 202651 -204
rect 202437 -294 202465 -266
rect 202499 -294 202527 -266
rect 202561 -294 202589 -266
rect 202623 -294 202651 -266
rect 204297 95147 204325 95175
rect 204359 95147 204387 95175
rect 204421 95147 204449 95175
rect 204483 95147 204511 95175
rect 204297 95085 204325 95113
rect 204359 95085 204387 95113
rect 204421 95085 204449 95113
rect 204483 95085 204511 95113
rect 204297 95023 204325 95051
rect 204359 95023 204387 95051
rect 204421 95023 204449 95051
rect 204483 95023 204511 95051
rect 204297 94961 204325 94989
rect 204359 94961 204387 94989
rect 204421 94961 204449 94989
rect 204483 94961 204511 94989
rect 204297 86147 204325 86175
rect 204359 86147 204387 86175
rect 204421 86147 204449 86175
rect 204483 86147 204511 86175
rect 204297 86085 204325 86113
rect 204359 86085 204387 86113
rect 204421 86085 204449 86113
rect 204483 86085 204511 86113
rect 204297 86023 204325 86051
rect 204359 86023 204387 86051
rect 204421 86023 204449 86051
rect 204483 86023 204511 86051
rect 204297 85961 204325 85989
rect 204359 85961 204387 85989
rect 204421 85961 204449 85989
rect 204483 85961 204511 85989
rect 204297 77147 204325 77175
rect 204359 77147 204387 77175
rect 204421 77147 204449 77175
rect 204483 77147 204511 77175
rect 204297 77085 204325 77113
rect 204359 77085 204387 77113
rect 204421 77085 204449 77113
rect 204483 77085 204511 77113
rect 204297 77023 204325 77051
rect 204359 77023 204387 77051
rect 204421 77023 204449 77051
rect 204483 77023 204511 77051
rect 204297 76961 204325 76989
rect 204359 76961 204387 76989
rect 204421 76961 204449 76989
rect 204483 76961 204511 76989
rect 204297 68147 204325 68175
rect 204359 68147 204387 68175
rect 204421 68147 204449 68175
rect 204483 68147 204511 68175
rect 204297 68085 204325 68113
rect 204359 68085 204387 68113
rect 204421 68085 204449 68113
rect 204483 68085 204511 68113
rect 204297 68023 204325 68051
rect 204359 68023 204387 68051
rect 204421 68023 204449 68051
rect 204483 68023 204511 68051
rect 204297 67961 204325 67989
rect 204359 67961 204387 67989
rect 204421 67961 204449 67989
rect 204483 67961 204511 67989
rect 204297 59147 204325 59175
rect 204359 59147 204387 59175
rect 204421 59147 204449 59175
rect 204483 59147 204511 59175
rect 204297 59085 204325 59113
rect 204359 59085 204387 59113
rect 204421 59085 204449 59113
rect 204483 59085 204511 59113
rect 204297 59023 204325 59051
rect 204359 59023 204387 59051
rect 204421 59023 204449 59051
rect 204483 59023 204511 59051
rect 204297 58961 204325 58989
rect 204359 58961 204387 58989
rect 204421 58961 204449 58989
rect 204483 58961 204511 58989
rect 204297 50147 204325 50175
rect 204359 50147 204387 50175
rect 204421 50147 204449 50175
rect 204483 50147 204511 50175
rect 204297 50085 204325 50113
rect 204359 50085 204387 50113
rect 204421 50085 204449 50113
rect 204483 50085 204511 50113
rect 204297 50023 204325 50051
rect 204359 50023 204387 50051
rect 204421 50023 204449 50051
rect 204483 50023 204511 50051
rect 204297 49961 204325 49989
rect 204359 49961 204387 49989
rect 204421 49961 204449 49989
rect 204483 49961 204511 49989
rect 204297 41147 204325 41175
rect 204359 41147 204387 41175
rect 204421 41147 204449 41175
rect 204483 41147 204511 41175
rect 204297 41085 204325 41113
rect 204359 41085 204387 41113
rect 204421 41085 204449 41113
rect 204483 41085 204511 41113
rect 204297 41023 204325 41051
rect 204359 41023 204387 41051
rect 204421 41023 204449 41051
rect 204483 41023 204511 41051
rect 204297 40961 204325 40989
rect 204359 40961 204387 40989
rect 204421 40961 204449 40989
rect 204483 40961 204511 40989
rect 204297 32147 204325 32175
rect 204359 32147 204387 32175
rect 204421 32147 204449 32175
rect 204483 32147 204511 32175
rect 204297 32085 204325 32113
rect 204359 32085 204387 32113
rect 204421 32085 204449 32113
rect 204483 32085 204511 32113
rect 204297 32023 204325 32051
rect 204359 32023 204387 32051
rect 204421 32023 204449 32051
rect 204483 32023 204511 32051
rect 204297 31961 204325 31989
rect 204359 31961 204387 31989
rect 204421 31961 204449 31989
rect 204483 31961 204511 31989
rect 204297 23147 204325 23175
rect 204359 23147 204387 23175
rect 204421 23147 204449 23175
rect 204483 23147 204511 23175
rect 204297 23085 204325 23113
rect 204359 23085 204387 23113
rect 204421 23085 204449 23113
rect 204483 23085 204511 23113
rect 204297 23023 204325 23051
rect 204359 23023 204387 23051
rect 204421 23023 204449 23051
rect 204483 23023 204511 23051
rect 204297 22961 204325 22989
rect 204359 22961 204387 22989
rect 204421 22961 204449 22989
rect 204483 22961 204511 22989
rect 204297 14147 204325 14175
rect 204359 14147 204387 14175
rect 204421 14147 204449 14175
rect 204483 14147 204511 14175
rect 204297 14085 204325 14113
rect 204359 14085 204387 14113
rect 204421 14085 204449 14113
rect 204483 14085 204511 14113
rect 204297 14023 204325 14051
rect 204359 14023 204387 14051
rect 204421 14023 204449 14051
rect 204483 14023 204511 14051
rect 204297 13961 204325 13989
rect 204359 13961 204387 13989
rect 204421 13961 204449 13989
rect 204483 13961 204511 13989
rect 204297 5147 204325 5175
rect 204359 5147 204387 5175
rect 204421 5147 204449 5175
rect 204483 5147 204511 5175
rect 204297 5085 204325 5113
rect 204359 5085 204387 5113
rect 204421 5085 204449 5113
rect 204483 5085 204511 5113
rect 204297 5023 204325 5051
rect 204359 5023 204387 5051
rect 204421 5023 204449 5051
rect 204483 5023 204511 5051
rect 204297 4961 204325 4989
rect 204359 4961 204387 4989
rect 204421 4961 204449 4989
rect 204483 4961 204511 4989
rect 204297 -588 204325 -560
rect 204359 -588 204387 -560
rect 204421 -588 204449 -560
rect 204483 -588 204511 -560
rect 204297 -650 204325 -622
rect 204359 -650 204387 -622
rect 204421 -650 204449 -622
rect 204483 -650 204511 -622
rect 204297 -712 204325 -684
rect 204359 -712 204387 -684
rect 204421 -712 204449 -684
rect 204483 -712 204511 -684
rect 204297 -774 204325 -746
rect 204359 -774 204387 -746
rect 204421 -774 204449 -746
rect 204483 -774 204511 -746
rect 217797 92147 217825 92175
rect 217859 92147 217887 92175
rect 217921 92147 217949 92175
rect 217983 92147 218011 92175
rect 217797 92085 217825 92113
rect 217859 92085 217887 92113
rect 217921 92085 217949 92113
rect 217983 92085 218011 92113
rect 217797 92023 217825 92051
rect 217859 92023 217887 92051
rect 217921 92023 217949 92051
rect 217983 92023 218011 92051
rect 217797 91961 217825 91989
rect 217859 91961 217887 91989
rect 217921 91961 217949 91989
rect 217983 91961 218011 91989
rect 217797 83147 217825 83175
rect 217859 83147 217887 83175
rect 217921 83147 217949 83175
rect 217983 83147 218011 83175
rect 217797 83085 217825 83113
rect 217859 83085 217887 83113
rect 217921 83085 217949 83113
rect 217983 83085 218011 83113
rect 217797 83023 217825 83051
rect 217859 83023 217887 83051
rect 217921 83023 217949 83051
rect 217983 83023 218011 83051
rect 217797 82961 217825 82989
rect 217859 82961 217887 82989
rect 217921 82961 217949 82989
rect 217983 82961 218011 82989
rect 217797 74147 217825 74175
rect 217859 74147 217887 74175
rect 217921 74147 217949 74175
rect 217983 74147 218011 74175
rect 217797 74085 217825 74113
rect 217859 74085 217887 74113
rect 217921 74085 217949 74113
rect 217983 74085 218011 74113
rect 217797 74023 217825 74051
rect 217859 74023 217887 74051
rect 217921 74023 217949 74051
rect 217983 74023 218011 74051
rect 217797 73961 217825 73989
rect 217859 73961 217887 73989
rect 217921 73961 217949 73989
rect 217983 73961 218011 73989
rect 217797 65147 217825 65175
rect 217859 65147 217887 65175
rect 217921 65147 217949 65175
rect 217983 65147 218011 65175
rect 217797 65085 217825 65113
rect 217859 65085 217887 65113
rect 217921 65085 217949 65113
rect 217983 65085 218011 65113
rect 217797 65023 217825 65051
rect 217859 65023 217887 65051
rect 217921 65023 217949 65051
rect 217983 65023 218011 65051
rect 217797 64961 217825 64989
rect 217859 64961 217887 64989
rect 217921 64961 217949 64989
rect 217983 64961 218011 64989
rect 217797 56147 217825 56175
rect 217859 56147 217887 56175
rect 217921 56147 217949 56175
rect 217983 56147 218011 56175
rect 217797 56085 217825 56113
rect 217859 56085 217887 56113
rect 217921 56085 217949 56113
rect 217983 56085 218011 56113
rect 217797 56023 217825 56051
rect 217859 56023 217887 56051
rect 217921 56023 217949 56051
rect 217983 56023 218011 56051
rect 217797 55961 217825 55989
rect 217859 55961 217887 55989
rect 217921 55961 217949 55989
rect 217983 55961 218011 55989
rect 217797 47147 217825 47175
rect 217859 47147 217887 47175
rect 217921 47147 217949 47175
rect 217983 47147 218011 47175
rect 217797 47085 217825 47113
rect 217859 47085 217887 47113
rect 217921 47085 217949 47113
rect 217983 47085 218011 47113
rect 217797 47023 217825 47051
rect 217859 47023 217887 47051
rect 217921 47023 217949 47051
rect 217983 47023 218011 47051
rect 217797 46961 217825 46989
rect 217859 46961 217887 46989
rect 217921 46961 217949 46989
rect 217983 46961 218011 46989
rect 217797 38147 217825 38175
rect 217859 38147 217887 38175
rect 217921 38147 217949 38175
rect 217983 38147 218011 38175
rect 217797 38085 217825 38113
rect 217859 38085 217887 38113
rect 217921 38085 217949 38113
rect 217983 38085 218011 38113
rect 217797 38023 217825 38051
rect 217859 38023 217887 38051
rect 217921 38023 217949 38051
rect 217983 38023 218011 38051
rect 217797 37961 217825 37989
rect 217859 37961 217887 37989
rect 217921 37961 217949 37989
rect 217983 37961 218011 37989
rect 217797 29147 217825 29175
rect 217859 29147 217887 29175
rect 217921 29147 217949 29175
rect 217983 29147 218011 29175
rect 217797 29085 217825 29113
rect 217859 29085 217887 29113
rect 217921 29085 217949 29113
rect 217983 29085 218011 29113
rect 217797 29023 217825 29051
rect 217859 29023 217887 29051
rect 217921 29023 217949 29051
rect 217983 29023 218011 29051
rect 217797 28961 217825 28989
rect 217859 28961 217887 28989
rect 217921 28961 217949 28989
rect 217983 28961 218011 28989
rect 217797 20147 217825 20175
rect 217859 20147 217887 20175
rect 217921 20147 217949 20175
rect 217983 20147 218011 20175
rect 217797 20085 217825 20113
rect 217859 20085 217887 20113
rect 217921 20085 217949 20113
rect 217983 20085 218011 20113
rect 217797 20023 217825 20051
rect 217859 20023 217887 20051
rect 217921 20023 217949 20051
rect 217983 20023 218011 20051
rect 217797 19961 217825 19989
rect 217859 19961 217887 19989
rect 217921 19961 217949 19989
rect 217983 19961 218011 19989
rect 217797 11147 217825 11175
rect 217859 11147 217887 11175
rect 217921 11147 217949 11175
rect 217983 11147 218011 11175
rect 217797 11085 217825 11113
rect 217859 11085 217887 11113
rect 217921 11085 217949 11113
rect 217983 11085 218011 11113
rect 217797 11023 217825 11051
rect 217859 11023 217887 11051
rect 217921 11023 217949 11051
rect 217983 11023 218011 11051
rect 217797 10961 217825 10989
rect 217859 10961 217887 10989
rect 217921 10961 217949 10989
rect 217983 10961 218011 10989
rect 217797 2147 217825 2175
rect 217859 2147 217887 2175
rect 217921 2147 217949 2175
rect 217983 2147 218011 2175
rect 217797 2085 217825 2113
rect 217859 2085 217887 2113
rect 217921 2085 217949 2113
rect 217983 2085 218011 2113
rect 217797 2023 217825 2051
rect 217859 2023 217887 2051
rect 217921 2023 217949 2051
rect 217983 2023 218011 2051
rect 217797 1961 217825 1989
rect 217859 1961 217887 1989
rect 217921 1961 217949 1989
rect 217983 1961 218011 1989
rect 217797 -108 217825 -80
rect 217859 -108 217887 -80
rect 217921 -108 217949 -80
rect 217983 -108 218011 -80
rect 217797 -170 217825 -142
rect 217859 -170 217887 -142
rect 217921 -170 217949 -142
rect 217983 -170 218011 -142
rect 217797 -232 217825 -204
rect 217859 -232 217887 -204
rect 217921 -232 217949 -204
rect 217983 -232 218011 -204
rect 217797 -294 217825 -266
rect 217859 -294 217887 -266
rect 217921 -294 217949 -266
rect 217983 -294 218011 -266
rect 219657 95147 219685 95175
rect 219719 95147 219747 95175
rect 219781 95147 219809 95175
rect 219843 95147 219871 95175
rect 219657 95085 219685 95113
rect 219719 95085 219747 95113
rect 219781 95085 219809 95113
rect 219843 95085 219871 95113
rect 219657 95023 219685 95051
rect 219719 95023 219747 95051
rect 219781 95023 219809 95051
rect 219843 95023 219871 95051
rect 219657 94961 219685 94989
rect 219719 94961 219747 94989
rect 219781 94961 219809 94989
rect 219843 94961 219871 94989
rect 219657 86147 219685 86175
rect 219719 86147 219747 86175
rect 219781 86147 219809 86175
rect 219843 86147 219871 86175
rect 219657 86085 219685 86113
rect 219719 86085 219747 86113
rect 219781 86085 219809 86113
rect 219843 86085 219871 86113
rect 219657 86023 219685 86051
rect 219719 86023 219747 86051
rect 219781 86023 219809 86051
rect 219843 86023 219871 86051
rect 219657 85961 219685 85989
rect 219719 85961 219747 85989
rect 219781 85961 219809 85989
rect 219843 85961 219871 85989
rect 219657 77147 219685 77175
rect 219719 77147 219747 77175
rect 219781 77147 219809 77175
rect 219843 77147 219871 77175
rect 219657 77085 219685 77113
rect 219719 77085 219747 77113
rect 219781 77085 219809 77113
rect 219843 77085 219871 77113
rect 219657 77023 219685 77051
rect 219719 77023 219747 77051
rect 219781 77023 219809 77051
rect 219843 77023 219871 77051
rect 219657 76961 219685 76989
rect 219719 76961 219747 76989
rect 219781 76961 219809 76989
rect 219843 76961 219871 76989
rect 219657 68147 219685 68175
rect 219719 68147 219747 68175
rect 219781 68147 219809 68175
rect 219843 68147 219871 68175
rect 219657 68085 219685 68113
rect 219719 68085 219747 68113
rect 219781 68085 219809 68113
rect 219843 68085 219871 68113
rect 219657 68023 219685 68051
rect 219719 68023 219747 68051
rect 219781 68023 219809 68051
rect 219843 68023 219871 68051
rect 219657 67961 219685 67989
rect 219719 67961 219747 67989
rect 219781 67961 219809 67989
rect 219843 67961 219871 67989
rect 219657 59147 219685 59175
rect 219719 59147 219747 59175
rect 219781 59147 219809 59175
rect 219843 59147 219871 59175
rect 219657 59085 219685 59113
rect 219719 59085 219747 59113
rect 219781 59085 219809 59113
rect 219843 59085 219871 59113
rect 219657 59023 219685 59051
rect 219719 59023 219747 59051
rect 219781 59023 219809 59051
rect 219843 59023 219871 59051
rect 219657 58961 219685 58989
rect 219719 58961 219747 58989
rect 219781 58961 219809 58989
rect 219843 58961 219871 58989
rect 219657 50147 219685 50175
rect 219719 50147 219747 50175
rect 219781 50147 219809 50175
rect 219843 50147 219871 50175
rect 219657 50085 219685 50113
rect 219719 50085 219747 50113
rect 219781 50085 219809 50113
rect 219843 50085 219871 50113
rect 219657 50023 219685 50051
rect 219719 50023 219747 50051
rect 219781 50023 219809 50051
rect 219843 50023 219871 50051
rect 219657 49961 219685 49989
rect 219719 49961 219747 49989
rect 219781 49961 219809 49989
rect 219843 49961 219871 49989
rect 219657 41147 219685 41175
rect 219719 41147 219747 41175
rect 219781 41147 219809 41175
rect 219843 41147 219871 41175
rect 219657 41085 219685 41113
rect 219719 41085 219747 41113
rect 219781 41085 219809 41113
rect 219843 41085 219871 41113
rect 219657 41023 219685 41051
rect 219719 41023 219747 41051
rect 219781 41023 219809 41051
rect 219843 41023 219871 41051
rect 219657 40961 219685 40989
rect 219719 40961 219747 40989
rect 219781 40961 219809 40989
rect 219843 40961 219871 40989
rect 219657 32147 219685 32175
rect 219719 32147 219747 32175
rect 219781 32147 219809 32175
rect 219843 32147 219871 32175
rect 219657 32085 219685 32113
rect 219719 32085 219747 32113
rect 219781 32085 219809 32113
rect 219843 32085 219871 32113
rect 219657 32023 219685 32051
rect 219719 32023 219747 32051
rect 219781 32023 219809 32051
rect 219843 32023 219871 32051
rect 219657 31961 219685 31989
rect 219719 31961 219747 31989
rect 219781 31961 219809 31989
rect 219843 31961 219871 31989
rect 219657 23147 219685 23175
rect 219719 23147 219747 23175
rect 219781 23147 219809 23175
rect 219843 23147 219871 23175
rect 219657 23085 219685 23113
rect 219719 23085 219747 23113
rect 219781 23085 219809 23113
rect 219843 23085 219871 23113
rect 219657 23023 219685 23051
rect 219719 23023 219747 23051
rect 219781 23023 219809 23051
rect 219843 23023 219871 23051
rect 219657 22961 219685 22989
rect 219719 22961 219747 22989
rect 219781 22961 219809 22989
rect 219843 22961 219871 22989
rect 219657 14147 219685 14175
rect 219719 14147 219747 14175
rect 219781 14147 219809 14175
rect 219843 14147 219871 14175
rect 219657 14085 219685 14113
rect 219719 14085 219747 14113
rect 219781 14085 219809 14113
rect 219843 14085 219871 14113
rect 219657 14023 219685 14051
rect 219719 14023 219747 14051
rect 219781 14023 219809 14051
rect 219843 14023 219871 14051
rect 219657 13961 219685 13989
rect 219719 13961 219747 13989
rect 219781 13961 219809 13989
rect 219843 13961 219871 13989
rect 219657 5147 219685 5175
rect 219719 5147 219747 5175
rect 219781 5147 219809 5175
rect 219843 5147 219871 5175
rect 219657 5085 219685 5113
rect 219719 5085 219747 5113
rect 219781 5085 219809 5113
rect 219843 5085 219871 5113
rect 219657 5023 219685 5051
rect 219719 5023 219747 5051
rect 219781 5023 219809 5051
rect 219843 5023 219871 5051
rect 219657 4961 219685 4989
rect 219719 4961 219747 4989
rect 219781 4961 219809 4989
rect 219843 4961 219871 4989
rect 219657 -588 219685 -560
rect 219719 -588 219747 -560
rect 219781 -588 219809 -560
rect 219843 -588 219871 -560
rect 219657 -650 219685 -622
rect 219719 -650 219747 -622
rect 219781 -650 219809 -622
rect 219843 -650 219871 -622
rect 219657 -712 219685 -684
rect 219719 -712 219747 -684
rect 219781 -712 219809 -684
rect 219843 -712 219871 -684
rect 219657 -774 219685 -746
rect 219719 -774 219747 -746
rect 219781 -774 219809 -746
rect 219843 -774 219871 -746
rect 233157 92147 233185 92175
rect 233219 92147 233247 92175
rect 233281 92147 233309 92175
rect 233343 92147 233371 92175
rect 233157 92085 233185 92113
rect 233219 92085 233247 92113
rect 233281 92085 233309 92113
rect 233343 92085 233371 92113
rect 233157 92023 233185 92051
rect 233219 92023 233247 92051
rect 233281 92023 233309 92051
rect 233343 92023 233371 92051
rect 233157 91961 233185 91989
rect 233219 91961 233247 91989
rect 233281 91961 233309 91989
rect 233343 91961 233371 91989
rect 233157 83147 233185 83175
rect 233219 83147 233247 83175
rect 233281 83147 233309 83175
rect 233343 83147 233371 83175
rect 233157 83085 233185 83113
rect 233219 83085 233247 83113
rect 233281 83085 233309 83113
rect 233343 83085 233371 83113
rect 233157 83023 233185 83051
rect 233219 83023 233247 83051
rect 233281 83023 233309 83051
rect 233343 83023 233371 83051
rect 233157 82961 233185 82989
rect 233219 82961 233247 82989
rect 233281 82961 233309 82989
rect 233343 82961 233371 82989
rect 233157 74147 233185 74175
rect 233219 74147 233247 74175
rect 233281 74147 233309 74175
rect 233343 74147 233371 74175
rect 233157 74085 233185 74113
rect 233219 74085 233247 74113
rect 233281 74085 233309 74113
rect 233343 74085 233371 74113
rect 233157 74023 233185 74051
rect 233219 74023 233247 74051
rect 233281 74023 233309 74051
rect 233343 74023 233371 74051
rect 233157 73961 233185 73989
rect 233219 73961 233247 73989
rect 233281 73961 233309 73989
rect 233343 73961 233371 73989
rect 233157 65147 233185 65175
rect 233219 65147 233247 65175
rect 233281 65147 233309 65175
rect 233343 65147 233371 65175
rect 233157 65085 233185 65113
rect 233219 65085 233247 65113
rect 233281 65085 233309 65113
rect 233343 65085 233371 65113
rect 233157 65023 233185 65051
rect 233219 65023 233247 65051
rect 233281 65023 233309 65051
rect 233343 65023 233371 65051
rect 233157 64961 233185 64989
rect 233219 64961 233247 64989
rect 233281 64961 233309 64989
rect 233343 64961 233371 64989
rect 233157 56147 233185 56175
rect 233219 56147 233247 56175
rect 233281 56147 233309 56175
rect 233343 56147 233371 56175
rect 233157 56085 233185 56113
rect 233219 56085 233247 56113
rect 233281 56085 233309 56113
rect 233343 56085 233371 56113
rect 233157 56023 233185 56051
rect 233219 56023 233247 56051
rect 233281 56023 233309 56051
rect 233343 56023 233371 56051
rect 233157 55961 233185 55989
rect 233219 55961 233247 55989
rect 233281 55961 233309 55989
rect 233343 55961 233371 55989
rect 233157 47147 233185 47175
rect 233219 47147 233247 47175
rect 233281 47147 233309 47175
rect 233343 47147 233371 47175
rect 233157 47085 233185 47113
rect 233219 47085 233247 47113
rect 233281 47085 233309 47113
rect 233343 47085 233371 47113
rect 233157 47023 233185 47051
rect 233219 47023 233247 47051
rect 233281 47023 233309 47051
rect 233343 47023 233371 47051
rect 233157 46961 233185 46989
rect 233219 46961 233247 46989
rect 233281 46961 233309 46989
rect 233343 46961 233371 46989
rect 233157 38147 233185 38175
rect 233219 38147 233247 38175
rect 233281 38147 233309 38175
rect 233343 38147 233371 38175
rect 233157 38085 233185 38113
rect 233219 38085 233247 38113
rect 233281 38085 233309 38113
rect 233343 38085 233371 38113
rect 233157 38023 233185 38051
rect 233219 38023 233247 38051
rect 233281 38023 233309 38051
rect 233343 38023 233371 38051
rect 233157 37961 233185 37989
rect 233219 37961 233247 37989
rect 233281 37961 233309 37989
rect 233343 37961 233371 37989
rect 233157 29147 233185 29175
rect 233219 29147 233247 29175
rect 233281 29147 233309 29175
rect 233343 29147 233371 29175
rect 233157 29085 233185 29113
rect 233219 29085 233247 29113
rect 233281 29085 233309 29113
rect 233343 29085 233371 29113
rect 233157 29023 233185 29051
rect 233219 29023 233247 29051
rect 233281 29023 233309 29051
rect 233343 29023 233371 29051
rect 233157 28961 233185 28989
rect 233219 28961 233247 28989
rect 233281 28961 233309 28989
rect 233343 28961 233371 28989
rect 233157 20147 233185 20175
rect 233219 20147 233247 20175
rect 233281 20147 233309 20175
rect 233343 20147 233371 20175
rect 233157 20085 233185 20113
rect 233219 20085 233247 20113
rect 233281 20085 233309 20113
rect 233343 20085 233371 20113
rect 233157 20023 233185 20051
rect 233219 20023 233247 20051
rect 233281 20023 233309 20051
rect 233343 20023 233371 20051
rect 233157 19961 233185 19989
rect 233219 19961 233247 19989
rect 233281 19961 233309 19989
rect 233343 19961 233371 19989
rect 233157 11147 233185 11175
rect 233219 11147 233247 11175
rect 233281 11147 233309 11175
rect 233343 11147 233371 11175
rect 233157 11085 233185 11113
rect 233219 11085 233247 11113
rect 233281 11085 233309 11113
rect 233343 11085 233371 11113
rect 233157 11023 233185 11051
rect 233219 11023 233247 11051
rect 233281 11023 233309 11051
rect 233343 11023 233371 11051
rect 233157 10961 233185 10989
rect 233219 10961 233247 10989
rect 233281 10961 233309 10989
rect 233343 10961 233371 10989
rect 233157 2147 233185 2175
rect 233219 2147 233247 2175
rect 233281 2147 233309 2175
rect 233343 2147 233371 2175
rect 233157 2085 233185 2113
rect 233219 2085 233247 2113
rect 233281 2085 233309 2113
rect 233343 2085 233371 2113
rect 233157 2023 233185 2051
rect 233219 2023 233247 2051
rect 233281 2023 233309 2051
rect 233343 2023 233371 2051
rect 233157 1961 233185 1989
rect 233219 1961 233247 1989
rect 233281 1961 233309 1989
rect 233343 1961 233371 1989
rect 233157 -108 233185 -80
rect 233219 -108 233247 -80
rect 233281 -108 233309 -80
rect 233343 -108 233371 -80
rect 233157 -170 233185 -142
rect 233219 -170 233247 -142
rect 233281 -170 233309 -142
rect 233343 -170 233371 -142
rect 233157 -232 233185 -204
rect 233219 -232 233247 -204
rect 233281 -232 233309 -204
rect 233343 -232 233371 -204
rect 233157 -294 233185 -266
rect 233219 -294 233247 -266
rect 233281 -294 233309 -266
rect 233343 -294 233371 -266
rect 235017 95147 235045 95175
rect 235079 95147 235107 95175
rect 235141 95147 235169 95175
rect 235203 95147 235231 95175
rect 235017 95085 235045 95113
rect 235079 95085 235107 95113
rect 235141 95085 235169 95113
rect 235203 95085 235231 95113
rect 235017 95023 235045 95051
rect 235079 95023 235107 95051
rect 235141 95023 235169 95051
rect 235203 95023 235231 95051
rect 235017 94961 235045 94989
rect 235079 94961 235107 94989
rect 235141 94961 235169 94989
rect 235203 94961 235231 94989
rect 235017 86147 235045 86175
rect 235079 86147 235107 86175
rect 235141 86147 235169 86175
rect 235203 86147 235231 86175
rect 235017 86085 235045 86113
rect 235079 86085 235107 86113
rect 235141 86085 235169 86113
rect 235203 86085 235231 86113
rect 235017 86023 235045 86051
rect 235079 86023 235107 86051
rect 235141 86023 235169 86051
rect 235203 86023 235231 86051
rect 235017 85961 235045 85989
rect 235079 85961 235107 85989
rect 235141 85961 235169 85989
rect 235203 85961 235231 85989
rect 235017 77147 235045 77175
rect 235079 77147 235107 77175
rect 235141 77147 235169 77175
rect 235203 77147 235231 77175
rect 235017 77085 235045 77113
rect 235079 77085 235107 77113
rect 235141 77085 235169 77113
rect 235203 77085 235231 77113
rect 235017 77023 235045 77051
rect 235079 77023 235107 77051
rect 235141 77023 235169 77051
rect 235203 77023 235231 77051
rect 235017 76961 235045 76989
rect 235079 76961 235107 76989
rect 235141 76961 235169 76989
rect 235203 76961 235231 76989
rect 235017 68147 235045 68175
rect 235079 68147 235107 68175
rect 235141 68147 235169 68175
rect 235203 68147 235231 68175
rect 235017 68085 235045 68113
rect 235079 68085 235107 68113
rect 235141 68085 235169 68113
rect 235203 68085 235231 68113
rect 235017 68023 235045 68051
rect 235079 68023 235107 68051
rect 235141 68023 235169 68051
rect 235203 68023 235231 68051
rect 235017 67961 235045 67989
rect 235079 67961 235107 67989
rect 235141 67961 235169 67989
rect 235203 67961 235231 67989
rect 235017 59147 235045 59175
rect 235079 59147 235107 59175
rect 235141 59147 235169 59175
rect 235203 59147 235231 59175
rect 235017 59085 235045 59113
rect 235079 59085 235107 59113
rect 235141 59085 235169 59113
rect 235203 59085 235231 59113
rect 235017 59023 235045 59051
rect 235079 59023 235107 59051
rect 235141 59023 235169 59051
rect 235203 59023 235231 59051
rect 235017 58961 235045 58989
rect 235079 58961 235107 58989
rect 235141 58961 235169 58989
rect 235203 58961 235231 58989
rect 235017 50147 235045 50175
rect 235079 50147 235107 50175
rect 235141 50147 235169 50175
rect 235203 50147 235231 50175
rect 235017 50085 235045 50113
rect 235079 50085 235107 50113
rect 235141 50085 235169 50113
rect 235203 50085 235231 50113
rect 235017 50023 235045 50051
rect 235079 50023 235107 50051
rect 235141 50023 235169 50051
rect 235203 50023 235231 50051
rect 235017 49961 235045 49989
rect 235079 49961 235107 49989
rect 235141 49961 235169 49989
rect 235203 49961 235231 49989
rect 235017 41147 235045 41175
rect 235079 41147 235107 41175
rect 235141 41147 235169 41175
rect 235203 41147 235231 41175
rect 235017 41085 235045 41113
rect 235079 41085 235107 41113
rect 235141 41085 235169 41113
rect 235203 41085 235231 41113
rect 235017 41023 235045 41051
rect 235079 41023 235107 41051
rect 235141 41023 235169 41051
rect 235203 41023 235231 41051
rect 235017 40961 235045 40989
rect 235079 40961 235107 40989
rect 235141 40961 235169 40989
rect 235203 40961 235231 40989
rect 235017 32147 235045 32175
rect 235079 32147 235107 32175
rect 235141 32147 235169 32175
rect 235203 32147 235231 32175
rect 235017 32085 235045 32113
rect 235079 32085 235107 32113
rect 235141 32085 235169 32113
rect 235203 32085 235231 32113
rect 235017 32023 235045 32051
rect 235079 32023 235107 32051
rect 235141 32023 235169 32051
rect 235203 32023 235231 32051
rect 235017 31961 235045 31989
rect 235079 31961 235107 31989
rect 235141 31961 235169 31989
rect 235203 31961 235231 31989
rect 235017 23147 235045 23175
rect 235079 23147 235107 23175
rect 235141 23147 235169 23175
rect 235203 23147 235231 23175
rect 235017 23085 235045 23113
rect 235079 23085 235107 23113
rect 235141 23085 235169 23113
rect 235203 23085 235231 23113
rect 235017 23023 235045 23051
rect 235079 23023 235107 23051
rect 235141 23023 235169 23051
rect 235203 23023 235231 23051
rect 235017 22961 235045 22989
rect 235079 22961 235107 22989
rect 235141 22961 235169 22989
rect 235203 22961 235231 22989
rect 235017 14147 235045 14175
rect 235079 14147 235107 14175
rect 235141 14147 235169 14175
rect 235203 14147 235231 14175
rect 235017 14085 235045 14113
rect 235079 14085 235107 14113
rect 235141 14085 235169 14113
rect 235203 14085 235231 14113
rect 235017 14023 235045 14051
rect 235079 14023 235107 14051
rect 235141 14023 235169 14051
rect 235203 14023 235231 14051
rect 235017 13961 235045 13989
rect 235079 13961 235107 13989
rect 235141 13961 235169 13989
rect 235203 13961 235231 13989
rect 235017 5147 235045 5175
rect 235079 5147 235107 5175
rect 235141 5147 235169 5175
rect 235203 5147 235231 5175
rect 235017 5085 235045 5113
rect 235079 5085 235107 5113
rect 235141 5085 235169 5113
rect 235203 5085 235231 5113
rect 235017 5023 235045 5051
rect 235079 5023 235107 5051
rect 235141 5023 235169 5051
rect 235203 5023 235231 5051
rect 235017 4961 235045 4989
rect 235079 4961 235107 4989
rect 235141 4961 235169 4989
rect 235203 4961 235231 4989
rect 235017 -588 235045 -560
rect 235079 -588 235107 -560
rect 235141 -588 235169 -560
rect 235203 -588 235231 -560
rect 235017 -650 235045 -622
rect 235079 -650 235107 -622
rect 235141 -650 235169 -622
rect 235203 -650 235231 -622
rect 235017 -712 235045 -684
rect 235079 -712 235107 -684
rect 235141 -712 235169 -684
rect 235203 -712 235231 -684
rect 235017 -774 235045 -746
rect 235079 -774 235107 -746
rect 235141 -774 235169 -746
rect 235203 -774 235231 -746
rect 248517 92147 248545 92175
rect 248579 92147 248607 92175
rect 248641 92147 248669 92175
rect 248703 92147 248731 92175
rect 248517 92085 248545 92113
rect 248579 92085 248607 92113
rect 248641 92085 248669 92113
rect 248703 92085 248731 92113
rect 248517 92023 248545 92051
rect 248579 92023 248607 92051
rect 248641 92023 248669 92051
rect 248703 92023 248731 92051
rect 248517 91961 248545 91989
rect 248579 91961 248607 91989
rect 248641 91961 248669 91989
rect 248703 91961 248731 91989
rect 248517 83147 248545 83175
rect 248579 83147 248607 83175
rect 248641 83147 248669 83175
rect 248703 83147 248731 83175
rect 248517 83085 248545 83113
rect 248579 83085 248607 83113
rect 248641 83085 248669 83113
rect 248703 83085 248731 83113
rect 248517 83023 248545 83051
rect 248579 83023 248607 83051
rect 248641 83023 248669 83051
rect 248703 83023 248731 83051
rect 248517 82961 248545 82989
rect 248579 82961 248607 82989
rect 248641 82961 248669 82989
rect 248703 82961 248731 82989
rect 248517 74147 248545 74175
rect 248579 74147 248607 74175
rect 248641 74147 248669 74175
rect 248703 74147 248731 74175
rect 248517 74085 248545 74113
rect 248579 74085 248607 74113
rect 248641 74085 248669 74113
rect 248703 74085 248731 74113
rect 248517 74023 248545 74051
rect 248579 74023 248607 74051
rect 248641 74023 248669 74051
rect 248703 74023 248731 74051
rect 248517 73961 248545 73989
rect 248579 73961 248607 73989
rect 248641 73961 248669 73989
rect 248703 73961 248731 73989
rect 248517 65147 248545 65175
rect 248579 65147 248607 65175
rect 248641 65147 248669 65175
rect 248703 65147 248731 65175
rect 248517 65085 248545 65113
rect 248579 65085 248607 65113
rect 248641 65085 248669 65113
rect 248703 65085 248731 65113
rect 248517 65023 248545 65051
rect 248579 65023 248607 65051
rect 248641 65023 248669 65051
rect 248703 65023 248731 65051
rect 248517 64961 248545 64989
rect 248579 64961 248607 64989
rect 248641 64961 248669 64989
rect 248703 64961 248731 64989
rect 248517 56147 248545 56175
rect 248579 56147 248607 56175
rect 248641 56147 248669 56175
rect 248703 56147 248731 56175
rect 248517 56085 248545 56113
rect 248579 56085 248607 56113
rect 248641 56085 248669 56113
rect 248703 56085 248731 56113
rect 248517 56023 248545 56051
rect 248579 56023 248607 56051
rect 248641 56023 248669 56051
rect 248703 56023 248731 56051
rect 248517 55961 248545 55989
rect 248579 55961 248607 55989
rect 248641 55961 248669 55989
rect 248703 55961 248731 55989
rect 248517 47147 248545 47175
rect 248579 47147 248607 47175
rect 248641 47147 248669 47175
rect 248703 47147 248731 47175
rect 248517 47085 248545 47113
rect 248579 47085 248607 47113
rect 248641 47085 248669 47113
rect 248703 47085 248731 47113
rect 248517 47023 248545 47051
rect 248579 47023 248607 47051
rect 248641 47023 248669 47051
rect 248703 47023 248731 47051
rect 248517 46961 248545 46989
rect 248579 46961 248607 46989
rect 248641 46961 248669 46989
rect 248703 46961 248731 46989
rect 248517 38147 248545 38175
rect 248579 38147 248607 38175
rect 248641 38147 248669 38175
rect 248703 38147 248731 38175
rect 248517 38085 248545 38113
rect 248579 38085 248607 38113
rect 248641 38085 248669 38113
rect 248703 38085 248731 38113
rect 248517 38023 248545 38051
rect 248579 38023 248607 38051
rect 248641 38023 248669 38051
rect 248703 38023 248731 38051
rect 248517 37961 248545 37989
rect 248579 37961 248607 37989
rect 248641 37961 248669 37989
rect 248703 37961 248731 37989
rect 248517 29147 248545 29175
rect 248579 29147 248607 29175
rect 248641 29147 248669 29175
rect 248703 29147 248731 29175
rect 248517 29085 248545 29113
rect 248579 29085 248607 29113
rect 248641 29085 248669 29113
rect 248703 29085 248731 29113
rect 248517 29023 248545 29051
rect 248579 29023 248607 29051
rect 248641 29023 248669 29051
rect 248703 29023 248731 29051
rect 248517 28961 248545 28989
rect 248579 28961 248607 28989
rect 248641 28961 248669 28989
rect 248703 28961 248731 28989
rect 248517 20147 248545 20175
rect 248579 20147 248607 20175
rect 248641 20147 248669 20175
rect 248703 20147 248731 20175
rect 248517 20085 248545 20113
rect 248579 20085 248607 20113
rect 248641 20085 248669 20113
rect 248703 20085 248731 20113
rect 248517 20023 248545 20051
rect 248579 20023 248607 20051
rect 248641 20023 248669 20051
rect 248703 20023 248731 20051
rect 248517 19961 248545 19989
rect 248579 19961 248607 19989
rect 248641 19961 248669 19989
rect 248703 19961 248731 19989
rect 248517 11147 248545 11175
rect 248579 11147 248607 11175
rect 248641 11147 248669 11175
rect 248703 11147 248731 11175
rect 248517 11085 248545 11113
rect 248579 11085 248607 11113
rect 248641 11085 248669 11113
rect 248703 11085 248731 11113
rect 248517 11023 248545 11051
rect 248579 11023 248607 11051
rect 248641 11023 248669 11051
rect 248703 11023 248731 11051
rect 248517 10961 248545 10989
rect 248579 10961 248607 10989
rect 248641 10961 248669 10989
rect 248703 10961 248731 10989
rect 248517 2147 248545 2175
rect 248579 2147 248607 2175
rect 248641 2147 248669 2175
rect 248703 2147 248731 2175
rect 248517 2085 248545 2113
rect 248579 2085 248607 2113
rect 248641 2085 248669 2113
rect 248703 2085 248731 2113
rect 248517 2023 248545 2051
rect 248579 2023 248607 2051
rect 248641 2023 248669 2051
rect 248703 2023 248731 2051
rect 248517 1961 248545 1989
rect 248579 1961 248607 1989
rect 248641 1961 248669 1989
rect 248703 1961 248731 1989
rect 248517 -108 248545 -80
rect 248579 -108 248607 -80
rect 248641 -108 248669 -80
rect 248703 -108 248731 -80
rect 248517 -170 248545 -142
rect 248579 -170 248607 -142
rect 248641 -170 248669 -142
rect 248703 -170 248731 -142
rect 248517 -232 248545 -204
rect 248579 -232 248607 -204
rect 248641 -232 248669 -204
rect 248703 -232 248731 -204
rect 248517 -294 248545 -266
rect 248579 -294 248607 -266
rect 248641 -294 248669 -266
rect 248703 -294 248731 -266
rect 250377 95147 250405 95175
rect 250439 95147 250467 95175
rect 250501 95147 250529 95175
rect 250563 95147 250591 95175
rect 250377 95085 250405 95113
rect 250439 95085 250467 95113
rect 250501 95085 250529 95113
rect 250563 95085 250591 95113
rect 250377 95023 250405 95051
rect 250439 95023 250467 95051
rect 250501 95023 250529 95051
rect 250563 95023 250591 95051
rect 250377 94961 250405 94989
rect 250439 94961 250467 94989
rect 250501 94961 250529 94989
rect 250563 94961 250591 94989
rect 250377 86147 250405 86175
rect 250439 86147 250467 86175
rect 250501 86147 250529 86175
rect 250563 86147 250591 86175
rect 250377 86085 250405 86113
rect 250439 86085 250467 86113
rect 250501 86085 250529 86113
rect 250563 86085 250591 86113
rect 250377 86023 250405 86051
rect 250439 86023 250467 86051
rect 250501 86023 250529 86051
rect 250563 86023 250591 86051
rect 250377 85961 250405 85989
rect 250439 85961 250467 85989
rect 250501 85961 250529 85989
rect 250563 85961 250591 85989
rect 250377 77147 250405 77175
rect 250439 77147 250467 77175
rect 250501 77147 250529 77175
rect 250563 77147 250591 77175
rect 250377 77085 250405 77113
rect 250439 77085 250467 77113
rect 250501 77085 250529 77113
rect 250563 77085 250591 77113
rect 250377 77023 250405 77051
rect 250439 77023 250467 77051
rect 250501 77023 250529 77051
rect 250563 77023 250591 77051
rect 250377 76961 250405 76989
rect 250439 76961 250467 76989
rect 250501 76961 250529 76989
rect 250563 76961 250591 76989
rect 250377 68147 250405 68175
rect 250439 68147 250467 68175
rect 250501 68147 250529 68175
rect 250563 68147 250591 68175
rect 250377 68085 250405 68113
rect 250439 68085 250467 68113
rect 250501 68085 250529 68113
rect 250563 68085 250591 68113
rect 250377 68023 250405 68051
rect 250439 68023 250467 68051
rect 250501 68023 250529 68051
rect 250563 68023 250591 68051
rect 250377 67961 250405 67989
rect 250439 67961 250467 67989
rect 250501 67961 250529 67989
rect 250563 67961 250591 67989
rect 250377 59147 250405 59175
rect 250439 59147 250467 59175
rect 250501 59147 250529 59175
rect 250563 59147 250591 59175
rect 250377 59085 250405 59113
rect 250439 59085 250467 59113
rect 250501 59085 250529 59113
rect 250563 59085 250591 59113
rect 250377 59023 250405 59051
rect 250439 59023 250467 59051
rect 250501 59023 250529 59051
rect 250563 59023 250591 59051
rect 250377 58961 250405 58989
rect 250439 58961 250467 58989
rect 250501 58961 250529 58989
rect 250563 58961 250591 58989
rect 250377 50147 250405 50175
rect 250439 50147 250467 50175
rect 250501 50147 250529 50175
rect 250563 50147 250591 50175
rect 250377 50085 250405 50113
rect 250439 50085 250467 50113
rect 250501 50085 250529 50113
rect 250563 50085 250591 50113
rect 250377 50023 250405 50051
rect 250439 50023 250467 50051
rect 250501 50023 250529 50051
rect 250563 50023 250591 50051
rect 250377 49961 250405 49989
rect 250439 49961 250467 49989
rect 250501 49961 250529 49989
rect 250563 49961 250591 49989
rect 250377 41147 250405 41175
rect 250439 41147 250467 41175
rect 250501 41147 250529 41175
rect 250563 41147 250591 41175
rect 250377 41085 250405 41113
rect 250439 41085 250467 41113
rect 250501 41085 250529 41113
rect 250563 41085 250591 41113
rect 250377 41023 250405 41051
rect 250439 41023 250467 41051
rect 250501 41023 250529 41051
rect 250563 41023 250591 41051
rect 250377 40961 250405 40989
rect 250439 40961 250467 40989
rect 250501 40961 250529 40989
rect 250563 40961 250591 40989
rect 250377 32147 250405 32175
rect 250439 32147 250467 32175
rect 250501 32147 250529 32175
rect 250563 32147 250591 32175
rect 250377 32085 250405 32113
rect 250439 32085 250467 32113
rect 250501 32085 250529 32113
rect 250563 32085 250591 32113
rect 250377 32023 250405 32051
rect 250439 32023 250467 32051
rect 250501 32023 250529 32051
rect 250563 32023 250591 32051
rect 250377 31961 250405 31989
rect 250439 31961 250467 31989
rect 250501 31961 250529 31989
rect 250563 31961 250591 31989
rect 250377 23147 250405 23175
rect 250439 23147 250467 23175
rect 250501 23147 250529 23175
rect 250563 23147 250591 23175
rect 250377 23085 250405 23113
rect 250439 23085 250467 23113
rect 250501 23085 250529 23113
rect 250563 23085 250591 23113
rect 250377 23023 250405 23051
rect 250439 23023 250467 23051
rect 250501 23023 250529 23051
rect 250563 23023 250591 23051
rect 250377 22961 250405 22989
rect 250439 22961 250467 22989
rect 250501 22961 250529 22989
rect 250563 22961 250591 22989
rect 250377 14147 250405 14175
rect 250439 14147 250467 14175
rect 250501 14147 250529 14175
rect 250563 14147 250591 14175
rect 250377 14085 250405 14113
rect 250439 14085 250467 14113
rect 250501 14085 250529 14113
rect 250563 14085 250591 14113
rect 250377 14023 250405 14051
rect 250439 14023 250467 14051
rect 250501 14023 250529 14051
rect 250563 14023 250591 14051
rect 250377 13961 250405 13989
rect 250439 13961 250467 13989
rect 250501 13961 250529 13989
rect 250563 13961 250591 13989
rect 250377 5147 250405 5175
rect 250439 5147 250467 5175
rect 250501 5147 250529 5175
rect 250563 5147 250591 5175
rect 250377 5085 250405 5113
rect 250439 5085 250467 5113
rect 250501 5085 250529 5113
rect 250563 5085 250591 5113
rect 250377 5023 250405 5051
rect 250439 5023 250467 5051
rect 250501 5023 250529 5051
rect 250563 5023 250591 5051
rect 250377 4961 250405 4989
rect 250439 4961 250467 4989
rect 250501 4961 250529 4989
rect 250563 4961 250591 4989
rect 250377 -588 250405 -560
rect 250439 -588 250467 -560
rect 250501 -588 250529 -560
rect 250563 -588 250591 -560
rect 250377 -650 250405 -622
rect 250439 -650 250467 -622
rect 250501 -650 250529 -622
rect 250563 -650 250591 -622
rect 250377 -712 250405 -684
rect 250439 -712 250467 -684
rect 250501 -712 250529 -684
rect 250563 -712 250591 -684
rect 250377 -774 250405 -746
rect 250439 -774 250467 -746
rect 250501 -774 250529 -746
rect 250563 -774 250591 -746
rect 263877 92147 263905 92175
rect 263939 92147 263967 92175
rect 264001 92147 264029 92175
rect 264063 92147 264091 92175
rect 263877 92085 263905 92113
rect 263939 92085 263967 92113
rect 264001 92085 264029 92113
rect 264063 92085 264091 92113
rect 263877 92023 263905 92051
rect 263939 92023 263967 92051
rect 264001 92023 264029 92051
rect 264063 92023 264091 92051
rect 263877 91961 263905 91989
rect 263939 91961 263967 91989
rect 264001 91961 264029 91989
rect 264063 91961 264091 91989
rect 263877 83147 263905 83175
rect 263939 83147 263967 83175
rect 264001 83147 264029 83175
rect 264063 83147 264091 83175
rect 263877 83085 263905 83113
rect 263939 83085 263967 83113
rect 264001 83085 264029 83113
rect 264063 83085 264091 83113
rect 263877 83023 263905 83051
rect 263939 83023 263967 83051
rect 264001 83023 264029 83051
rect 264063 83023 264091 83051
rect 263877 82961 263905 82989
rect 263939 82961 263967 82989
rect 264001 82961 264029 82989
rect 264063 82961 264091 82989
rect 263877 74147 263905 74175
rect 263939 74147 263967 74175
rect 264001 74147 264029 74175
rect 264063 74147 264091 74175
rect 263877 74085 263905 74113
rect 263939 74085 263967 74113
rect 264001 74085 264029 74113
rect 264063 74085 264091 74113
rect 263877 74023 263905 74051
rect 263939 74023 263967 74051
rect 264001 74023 264029 74051
rect 264063 74023 264091 74051
rect 263877 73961 263905 73989
rect 263939 73961 263967 73989
rect 264001 73961 264029 73989
rect 264063 73961 264091 73989
rect 263877 65147 263905 65175
rect 263939 65147 263967 65175
rect 264001 65147 264029 65175
rect 264063 65147 264091 65175
rect 263877 65085 263905 65113
rect 263939 65085 263967 65113
rect 264001 65085 264029 65113
rect 264063 65085 264091 65113
rect 263877 65023 263905 65051
rect 263939 65023 263967 65051
rect 264001 65023 264029 65051
rect 264063 65023 264091 65051
rect 263877 64961 263905 64989
rect 263939 64961 263967 64989
rect 264001 64961 264029 64989
rect 264063 64961 264091 64989
rect 263877 56147 263905 56175
rect 263939 56147 263967 56175
rect 264001 56147 264029 56175
rect 264063 56147 264091 56175
rect 263877 56085 263905 56113
rect 263939 56085 263967 56113
rect 264001 56085 264029 56113
rect 264063 56085 264091 56113
rect 263877 56023 263905 56051
rect 263939 56023 263967 56051
rect 264001 56023 264029 56051
rect 264063 56023 264091 56051
rect 263877 55961 263905 55989
rect 263939 55961 263967 55989
rect 264001 55961 264029 55989
rect 264063 55961 264091 55989
rect 263877 47147 263905 47175
rect 263939 47147 263967 47175
rect 264001 47147 264029 47175
rect 264063 47147 264091 47175
rect 263877 47085 263905 47113
rect 263939 47085 263967 47113
rect 264001 47085 264029 47113
rect 264063 47085 264091 47113
rect 263877 47023 263905 47051
rect 263939 47023 263967 47051
rect 264001 47023 264029 47051
rect 264063 47023 264091 47051
rect 263877 46961 263905 46989
rect 263939 46961 263967 46989
rect 264001 46961 264029 46989
rect 264063 46961 264091 46989
rect 263877 38147 263905 38175
rect 263939 38147 263967 38175
rect 264001 38147 264029 38175
rect 264063 38147 264091 38175
rect 263877 38085 263905 38113
rect 263939 38085 263967 38113
rect 264001 38085 264029 38113
rect 264063 38085 264091 38113
rect 263877 38023 263905 38051
rect 263939 38023 263967 38051
rect 264001 38023 264029 38051
rect 264063 38023 264091 38051
rect 263877 37961 263905 37989
rect 263939 37961 263967 37989
rect 264001 37961 264029 37989
rect 264063 37961 264091 37989
rect 263877 29147 263905 29175
rect 263939 29147 263967 29175
rect 264001 29147 264029 29175
rect 264063 29147 264091 29175
rect 263877 29085 263905 29113
rect 263939 29085 263967 29113
rect 264001 29085 264029 29113
rect 264063 29085 264091 29113
rect 263877 29023 263905 29051
rect 263939 29023 263967 29051
rect 264001 29023 264029 29051
rect 264063 29023 264091 29051
rect 263877 28961 263905 28989
rect 263939 28961 263967 28989
rect 264001 28961 264029 28989
rect 264063 28961 264091 28989
rect 263877 20147 263905 20175
rect 263939 20147 263967 20175
rect 264001 20147 264029 20175
rect 264063 20147 264091 20175
rect 263877 20085 263905 20113
rect 263939 20085 263967 20113
rect 264001 20085 264029 20113
rect 264063 20085 264091 20113
rect 263877 20023 263905 20051
rect 263939 20023 263967 20051
rect 264001 20023 264029 20051
rect 264063 20023 264091 20051
rect 263877 19961 263905 19989
rect 263939 19961 263967 19989
rect 264001 19961 264029 19989
rect 264063 19961 264091 19989
rect 263877 11147 263905 11175
rect 263939 11147 263967 11175
rect 264001 11147 264029 11175
rect 264063 11147 264091 11175
rect 263877 11085 263905 11113
rect 263939 11085 263967 11113
rect 264001 11085 264029 11113
rect 264063 11085 264091 11113
rect 263877 11023 263905 11051
rect 263939 11023 263967 11051
rect 264001 11023 264029 11051
rect 264063 11023 264091 11051
rect 263877 10961 263905 10989
rect 263939 10961 263967 10989
rect 264001 10961 264029 10989
rect 264063 10961 264091 10989
rect 263877 2147 263905 2175
rect 263939 2147 263967 2175
rect 264001 2147 264029 2175
rect 264063 2147 264091 2175
rect 263877 2085 263905 2113
rect 263939 2085 263967 2113
rect 264001 2085 264029 2113
rect 264063 2085 264091 2113
rect 263877 2023 263905 2051
rect 263939 2023 263967 2051
rect 264001 2023 264029 2051
rect 264063 2023 264091 2051
rect 263877 1961 263905 1989
rect 263939 1961 263967 1989
rect 264001 1961 264029 1989
rect 264063 1961 264091 1989
rect 263877 -108 263905 -80
rect 263939 -108 263967 -80
rect 264001 -108 264029 -80
rect 264063 -108 264091 -80
rect 263877 -170 263905 -142
rect 263939 -170 263967 -142
rect 264001 -170 264029 -142
rect 264063 -170 264091 -142
rect 263877 -232 263905 -204
rect 263939 -232 263967 -204
rect 264001 -232 264029 -204
rect 264063 -232 264091 -204
rect 263877 -294 263905 -266
rect 263939 -294 263967 -266
rect 264001 -294 264029 -266
rect 264063 -294 264091 -266
rect 265737 95147 265765 95175
rect 265799 95147 265827 95175
rect 265861 95147 265889 95175
rect 265923 95147 265951 95175
rect 265737 95085 265765 95113
rect 265799 95085 265827 95113
rect 265861 95085 265889 95113
rect 265923 95085 265951 95113
rect 265737 95023 265765 95051
rect 265799 95023 265827 95051
rect 265861 95023 265889 95051
rect 265923 95023 265951 95051
rect 265737 94961 265765 94989
rect 265799 94961 265827 94989
rect 265861 94961 265889 94989
rect 265923 94961 265951 94989
rect 265737 86147 265765 86175
rect 265799 86147 265827 86175
rect 265861 86147 265889 86175
rect 265923 86147 265951 86175
rect 265737 86085 265765 86113
rect 265799 86085 265827 86113
rect 265861 86085 265889 86113
rect 265923 86085 265951 86113
rect 265737 86023 265765 86051
rect 265799 86023 265827 86051
rect 265861 86023 265889 86051
rect 265923 86023 265951 86051
rect 265737 85961 265765 85989
rect 265799 85961 265827 85989
rect 265861 85961 265889 85989
rect 265923 85961 265951 85989
rect 265737 77147 265765 77175
rect 265799 77147 265827 77175
rect 265861 77147 265889 77175
rect 265923 77147 265951 77175
rect 265737 77085 265765 77113
rect 265799 77085 265827 77113
rect 265861 77085 265889 77113
rect 265923 77085 265951 77113
rect 265737 77023 265765 77051
rect 265799 77023 265827 77051
rect 265861 77023 265889 77051
rect 265923 77023 265951 77051
rect 265737 76961 265765 76989
rect 265799 76961 265827 76989
rect 265861 76961 265889 76989
rect 265923 76961 265951 76989
rect 265737 68147 265765 68175
rect 265799 68147 265827 68175
rect 265861 68147 265889 68175
rect 265923 68147 265951 68175
rect 265737 68085 265765 68113
rect 265799 68085 265827 68113
rect 265861 68085 265889 68113
rect 265923 68085 265951 68113
rect 265737 68023 265765 68051
rect 265799 68023 265827 68051
rect 265861 68023 265889 68051
rect 265923 68023 265951 68051
rect 265737 67961 265765 67989
rect 265799 67961 265827 67989
rect 265861 67961 265889 67989
rect 265923 67961 265951 67989
rect 265737 59147 265765 59175
rect 265799 59147 265827 59175
rect 265861 59147 265889 59175
rect 265923 59147 265951 59175
rect 265737 59085 265765 59113
rect 265799 59085 265827 59113
rect 265861 59085 265889 59113
rect 265923 59085 265951 59113
rect 265737 59023 265765 59051
rect 265799 59023 265827 59051
rect 265861 59023 265889 59051
rect 265923 59023 265951 59051
rect 265737 58961 265765 58989
rect 265799 58961 265827 58989
rect 265861 58961 265889 58989
rect 265923 58961 265951 58989
rect 265737 50147 265765 50175
rect 265799 50147 265827 50175
rect 265861 50147 265889 50175
rect 265923 50147 265951 50175
rect 265737 50085 265765 50113
rect 265799 50085 265827 50113
rect 265861 50085 265889 50113
rect 265923 50085 265951 50113
rect 265737 50023 265765 50051
rect 265799 50023 265827 50051
rect 265861 50023 265889 50051
rect 265923 50023 265951 50051
rect 265737 49961 265765 49989
rect 265799 49961 265827 49989
rect 265861 49961 265889 49989
rect 265923 49961 265951 49989
rect 265737 41147 265765 41175
rect 265799 41147 265827 41175
rect 265861 41147 265889 41175
rect 265923 41147 265951 41175
rect 265737 41085 265765 41113
rect 265799 41085 265827 41113
rect 265861 41085 265889 41113
rect 265923 41085 265951 41113
rect 265737 41023 265765 41051
rect 265799 41023 265827 41051
rect 265861 41023 265889 41051
rect 265923 41023 265951 41051
rect 265737 40961 265765 40989
rect 265799 40961 265827 40989
rect 265861 40961 265889 40989
rect 265923 40961 265951 40989
rect 265737 32147 265765 32175
rect 265799 32147 265827 32175
rect 265861 32147 265889 32175
rect 265923 32147 265951 32175
rect 265737 32085 265765 32113
rect 265799 32085 265827 32113
rect 265861 32085 265889 32113
rect 265923 32085 265951 32113
rect 265737 32023 265765 32051
rect 265799 32023 265827 32051
rect 265861 32023 265889 32051
rect 265923 32023 265951 32051
rect 265737 31961 265765 31989
rect 265799 31961 265827 31989
rect 265861 31961 265889 31989
rect 265923 31961 265951 31989
rect 265737 23147 265765 23175
rect 265799 23147 265827 23175
rect 265861 23147 265889 23175
rect 265923 23147 265951 23175
rect 265737 23085 265765 23113
rect 265799 23085 265827 23113
rect 265861 23085 265889 23113
rect 265923 23085 265951 23113
rect 265737 23023 265765 23051
rect 265799 23023 265827 23051
rect 265861 23023 265889 23051
rect 265923 23023 265951 23051
rect 265737 22961 265765 22989
rect 265799 22961 265827 22989
rect 265861 22961 265889 22989
rect 265923 22961 265951 22989
rect 265737 14147 265765 14175
rect 265799 14147 265827 14175
rect 265861 14147 265889 14175
rect 265923 14147 265951 14175
rect 265737 14085 265765 14113
rect 265799 14085 265827 14113
rect 265861 14085 265889 14113
rect 265923 14085 265951 14113
rect 265737 14023 265765 14051
rect 265799 14023 265827 14051
rect 265861 14023 265889 14051
rect 265923 14023 265951 14051
rect 265737 13961 265765 13989
rect 265799 13961 265827 13989
rect 265861 13961 265889 13989
rect 265923 13961 265951 13989
rect 265737 5147 265765 5175
rect 265799 5147 265827 5175
rect 265861 5147 265889 5175
rect 265923 5147 265951 5175
rect 265737 5085 265765 5113
rect 265799 5085 265827 5113
rect 265861 5085 265889 5113
rect 265923 5085 265951 5113
rect 265737 5023 265765 5051
rect 265799 5023 265827 5051
rect 265861 5023 265889 5051
rect 265923 5023 265951 5051
rect 265737 4961 265765 4989
rect 265799 4961 265827 4989
rect 265861 4961 265889 4989
rect 265923 4961 265951 4989
rect 265737 -588 265765 -560
rect 265799 -588 265827 -560
rect 265861 -588 265889 -560
rect 265923 -588 265951 -560
rect 265737 -650 265765 -622
rect 265799 -650 265827 -622
rect 265861 -650 265889 -622
rect 265923 -650 265951 -622
rect 265737 -712 265765 -684
rect 265799 -712 265827 -684
rect 265861 -712 265889 -684
rect 265923 -712 265951 -684
rect 265737 -774 265765 -746
rect 265799 -774 265827 -746
rect 265861 -774 265889 -746
rect 265923 -774 265951 -746
rect 279237 92147 279265 92175
rect 279299 92147 279327 92175
rect 279361 92147 279389 92175
rect 279423 92147 279451 92175
rect 279237 92085 279265 92113
rect 279299 92085 279327 92113
rect 279361 92085 279389 92113
rect 279423 92085 279451 92113
rect 279237 92023 279265 92051
rect 279299 92023 279327 92051
rect 279361 92023 279389 92051
rect 279423 92023 279451 92051
rect 279237 91961 279265 91989
rect 279299 91961 279327 91989
rect 279361 91961 279389 91989
rect 279423 91961 279451 91989
rect 279237 83147 279265 83175
rect 279299 83147 279327 83175
rect 279361 83147 279389 83175
rect 279423 83147 279451 83175
rect 279237 83085 279265 83113
rect 279299 83085 279327 83113
rect 279361 83085 279389 83113
rect 279423 83085 279451 83113
rect 279237 83023 279265 83051
rect 279299 83023 279327 83051
rect 279361 83023 279389 83051
rect 279423 83023 279451 83051
rect 279237 82961 279265 82989
rect 279299 82961 279327 82989
rect 279361 82961 279389 82989
rect 279423 82961 279451 82989
rect 279237 74147 279265 74175
rect 279299 74147 279327 74175
rect 279361 74147 279389 74175
rect 279423 74147 279451 74175
rect 279237 74085 279265 74113
rect 279299 74085 279327 74113
rect 279361 74085 279389 74113
rect 279423 74085 279451 74113
rect 279237 74023 279265 74051
rect 279299 74023 279327 74051
rect 279361 74023 279389 74051
rect 279423 74023 279451 74051
rect 279237 73961 279265 73989
rect 279299 73961 279327 73989
rect 279361 73961 279389 73989
rect 279423 73961 279451 73989
rect 279237 65147 279265 65175
rect 279299 65147 279327 65175
rect 279361 65147 279389 65175
rect 279423 65147 279451 65175
rect 279237 65085 279265 65113
rect 279299 65085 279327 65113
rect 279361 65085 279389 65113
rect 279423 65085 279451 65113
rect 279237 65023 279265 65051
rect 279299 65023 279327 65051
rect 279361 65023 279389 65051
rect 279423 65023 279451 65051
rect 279237 64961 279265 64989
rect 279299 64961 279327 64989
rect 279361 64961 279389 64989
rect 279423 64961 279451 64989
rect 279237 56147 279265 56175
rect 279299 56147 279327 56175
rect 279361 56147 279389 56175
rect 279423 56147 279451 56175
rect 279237 56085 279265 56113
rect 279299 56085 279327 56113
rect 279361 56085 279389 56113
rect 279423 56085 279451 56113
rect 279237 56023 279265 56051
rect 279299 56023 279327 56051
rect 279361 56023 279389 56051
rect 279423 56023 279451 56051
rect 279237 55961 279265 55989
rect 279299 55961 279327 55989
rect 279361 55961 279389 55989
rect 279423 55961 279451 55989
rect 279237 47147 279265 47175
rect 279299 47147 279327 47175
rect 279361 47147 279389 47175
rect 279423 47147 279451 47175
rect 279237 47085 279265 47113
rect 279299 47085 279327 47113
rect 279361 47085 279389 47113
rect 279423 47085 279451 47113
rect 279237 47023 279265 47051
rect 279299 47023 279327 47051
rect 279361 47023 279389 47051
rect 279423 47023 279451 47051
rect 279237 46961 279265 46989
rect 279299 46961 279327 46989
rect 279361 46961 279389 46989
rect 279423 46961 279451 46989
rect 279237 38147 279265 38175
rect 279299 38147 279327 38175
rect 279361 38147 279389 38175
rect 279423 38147 279451 38175
rect 279237 38085 279265 38113
rect 279299 38085 279327 38113
rect 279361 38085 279389 38113
rect 279423 38085 279451 38113
rect 279237 38023 279265 38051
rect 279299 38023 279327 38051
rect 279361 38023 279389 38051
rect 279423 38023 279451 38051
rect 279237 37961 279265 37989
rect 279299 37961 279327 37989
rect 279361 37961 279389 37989
rect 279423 37961 279451 37989
rect 279237 29147 279265 29175
rect 279299 29147 279327 29175
rect 279361 29147 279389 29175
rect 279423 29147 279451 29175
rect 279237 29085 279265 29113
rect 279299 29085 279327 29113
rect 279361 29085 279389 29113
rect 279423 29085 279451 29113
rect 279237 29023 279265 29051
rect 279299 29023 279327 29051
rect 279361 29023 279389 29051
rect 279423 29023 279451 29051
rect 279237 28961 279265 28989
rect 279299 28961 279327 28989
rect 279361 28961 279389 28989
rect 279423 28961 279451 28989
rect 279237 20147 279265 20175
rect 279299 20147 279327 20175
rect 279361 20147 279389 20175
rect 279423 20147 279451 20175
rect 279237 20085 279265 20113
rect 279299 20085 279327 20113
rect 279361 20085 279389 20113
rect 279423 20085 279451 20113
rect 279237 20023 279265 20051
rect 279299 20023 279327 20051
rect 279361 20023 279389 20051
rect 279423 20023 279451 20051
rect 279237 19961 279265 19989
rect 279299 19961 279327 19989
rect 279361 19961 279389 19989
rect 279423 19961 279451 19989
rect 279237 11147 279265 11175
rect 279299 11147 279327 11175
rect 279361 11147 279389 11175
rect 279423 11147 279451 11175
rect 279237 11085 279265 11113
rect 279299 11085 279327 11113
rect 279361 11085 279389 11113
rect 279423 11085 279451 11113
rect 279237 11023 279265 11051
rect 279299 11023 279327 11051
rect 279361 11023 279389 11051
rect 279423 11023 279451 11051
rect 279237 10961 279265 10989
rect 279299 10961 279327 10989
rect 279361 10961 279389 10989
rect 279423 10961 279451 10989
rect 279237 2147 279265 2175
rect 279299 2147 279327 2175
rect 279361 2147 279389 2175
rect 279423 2147 279451 2175
rect 279237 2085 279265 2113
rect 279299 2085 279327 2113
rect 279361 2085 279389 2113
rect 279423 2085 279451 2113
rect 279237 2023 279265 2051
rect 279299 2023 279327 2051
rect 279361 2023 279389 2051
rect 279423 2023 279451 2051
rect 279237 1961 279265 1989
rect 279299 1961 279327 1989
rect 279361 1961 279389 1989
rect 279423 1961 279451 1989
rect 279237 -108 279265 -80
rect 279299 -108 279327 -80
rect 279361 -108 279389 -80
rect 279423 -108 279451 -80
rect 279237 -170 279265 -142
rect 279299 -170 279327 -142
rect 279361 -170 279389 -142
rect 279423 -170 279451 -142
rect 279237 -232 279265 -204
rect 279299 -232 279327 -204
rect 279361 -232 279389 -204
rect 279423 -232 279451 -204
rect 279237 -294 279265 -266
rect 279299 -294 279327 -266
rect 279361 -294 279389 -266
rect 279423 -294 279451 -266
rect 281097 299058 281125 299086
rect 281159 299058 281187 299086
rect 281221 299058 281249 299086
rect 281283 299058 281311 299086
rect 281097 298996 281125 299024
rect 281159 298996 281187 299024
rect 281221 298996 281249 299024
rect 281283 298996 281311 299024
rect 281097 298934 281125 298962
rect 281159 298934 281187 298962
rect 281221 298934 281249 298962
rect 281283 298934 281311 298962
rect 281097 298872 281125 298900
rect 281159 298872 281187 298900
rect 281221 298872 281249 298900
rect 281283 298872 281311 298900
rect 281097 293147 281125 293175
rect 281159 293147 281187 293175
rect 281221 293147 281249 293175
rect 281283 293147 281311 293175
rect 281097 293085 281125 293113
rect 281159 293085 281187 293113
rect 281221 293085 281249 293113
rect 281283 293085 281311 293113
rect 281097 293023 281125 293051
rect 281159 293023 281187 293051
rect 281221 293023 281249 293051
rect 281283 293023 281311 293051
rect 281097 292961 281125 292989
rect 281159 292961 281187 292989
rect 281221 292961 281249 292989
rect 281283 292961 281311 292989
rect 281097 284147 281125 284175
rect 281159 284147 281187 284175
rect 281221 284147 281249 284175
rect 281283 284147 281311 284175
rect 281097 284085 281125 284113
rect 281159 284085 281187 284113
rect 281221 284085 281249 284113
rect 281283 284085 281311 284113
rect 281097 284023 281125 284051
rect 281159 284023 281187 284051
rect 281221 284023 281249 284051
rect 281283 284023 281311 284051
rect 281097 283961 281125 283989
rect 281159 283961 281187 283989
rect 281221 283961 281249 283989
rect 281283 283961 281311 283989
rect 281097 275147 281125 275175
rect 281159 275147 281187 275175
rect 281221 275147 281249 275175
rect 281283 275147 281311 275175
rect 281097 275085 281125 275113
rect 281159 275085 281187 275113
rect 281221 275085 281249 275113
rect 281283 275085 281311 275113
rect 281097 275023 281125 275051
rect 281159 275023 281187 275051
rect 281221 275023 281249 275051
rect 281283 275023 281311 275051
rect 294597 298578 294625 298606
rect 294659 298578 294687 298606
rect 294721 298578 294749 298606
rect 294783 298578 294811 298606
rect 294597 298516 294625 298544
rect 294659 298516 294687 298544
rect 294721 298516 294749 298544
rect 294783 298516 294811 298544
rect 294597 298454 294625 298482
rect 294659 298454 294687 298482
rect 294721 298454 294749 298482
rect 294783 298454 294811 298482
rect 294597 298392 294625 298420
rect 294659 298392 294687 298420
rect 294721 298392 294749 298420
rect 294783 298392 294811 298420
rect 294597 290147 294625 290175
rect 294659 290147 294687 290175
rect 294721 290147 294749 290175
rect 294783 290147 294811 290175
rect 294597 290085 294625 290113
rect 294659 290085 294687 290113
rect 294721 290085 294749 290113
rect 294783 290085 294811 290113
rect 294597 290023 294625 290051
rect 294659 290023 294687 290051
rect 294721 290023 294749 290051
rect 294783 290023 294811 290051
rect 294597 289961 294625 289989
rect 294659 289961 294687 289989
rect 294721 289961 294749 289989
rect 294783 289961 294811 289989
rect 294597 281147 294625 281175
rect 294659 281147 294687 281175
rect 294721 281147 294749 281175
rect 294783 281147 294811 281175
rect 294597 281085 294625 281113
rect 294659 281085 294687 281113
rect 294721 281085 294749 281113
rect 294783 281085 294811 281113
rect 294597 281023 294625 281051
rect 294659 281023 294687 281051
rect 294721 281023 294749 281051
rect 294783 281023 294811 281051
rect 294597 280961 294625 280989
rect 294659 280961 294687 280989
rect 294721 280961 294749 280989
rect 294783 280961 294811 280989
rect 281097 274961 281125 274989
rect 281159 274961 281187 274989
rect 281221 274961 281249 274989
rect 281283 274961 281311 274989
rect 281097 266147 281125 266175
rect 281159 266147 281187 266175
rect 281221 266147 281249 266175
rect 281283 266147 281311 266175
rect 281097 266085 281125 266113
rect 281159 266085 281187 266113
rect 281221 266085 281249 266113
rect 281283 266085 281311 266113
rect 281097 266023 281125 266051
rect 281159 266023 281187 266051
rect 281221 266023 281249 266051
rect 281283 266023 281311 266051
rect 281097 265961 281125 265989
rect 281159 265961 281187 265989
rect 281221 265961 281249 265989
rect 281283 265961 281311 265989
rect 281097 257147 281125 257175
rect 281159 257147 281187 257175
rect 281221 257147 281249 257175
rect 281283 257147 281311 257175
rect 281097 257085 281125 257113
rect 281159 257085 281187 257113
rect 281221 257085 281249 257113
rect 281283 257085 281311 257113
rect 281097 257023 281125 257051
rect 281159 257023 281187 257051
rect 281221 257023 281249 257051
rect 281283 257023 281311 257051
rect 281097 256961 281125 256989
rect 281159 256961 281187 256989
rect 281221 256961 281249 256989
rect 281283 256961 281311 256989
rect 281097 248147 281125 248175
rect 281159 248147 281187 248175
rect 281221 248147 281249 248175
rect 281283 248147 281311 248175
rect 281097 248085 281125 248113
rect 281159 248085 281187 248113
rect 281221 248085 281249 248113
rect 281283 248085 281311 248113
rect 281097 248023 281125 248051
rect 281159 248023 281187 248051
rect 281221 248023 281249 248051
rect 281283 248023 281311 248051
rect 281097 247961 281125 247989
rect 281159 247961 281187 247989
rect 281221 247961 281249 247989
rect 281283 247961 281311 247989
rect 281097 239147 281125 239175
rect 281159 239147 281187 239175
rect 281221 239147 281249 239175
rect 281283 239147 281311 239175
rect 281097 239085 281125 239113
rect 281159 239085 281187 239113
rect 281221 239085 281249 239113
rect 281283 239085 281311 239113
rect 281097 239023 281125 239051
rect 281159 239023 281187 239051
rect 281221 239023 281249 239051
rect 281283 239023 281311 239051
rect 281097 238961 281125 238989
rect 281159 238961 281187 238989
rect 281221 238961 281249 238989
rect 281283 238961 281311 238989
rect 281097 230147 281125 230175
rect 281159 230147 281187 230175
rect 281221 230147 281249 230175
rect 281283 230147 281311 230175
rect 281097 230085 281125 230113
rect 281159 230085 281187 230113
rect 281221 230085 281249 230113
rect 281283 230085 281311 230113
rect 281097 230023 281125 230051
rect 281159 230023 281187 230051
rect 281221 230023 281249 230051
rect 281283 230023 281311 230051
rect 281097 229961 281125 229989
rect 281159 229961 281187 229989
rect 281221 229961 281249 229989
rect 281283 229961 281311 229989
rect 281097 221147 281125 221175
rect 281159 221147 281187 221175
rect 281221 221147 281249 221175
rect 281283 221147 281311 221175
rect 281097 221085 281125 221113
rect 281159 221085 281187 221113
rect 281221 221085 281249 221113
rect 281283 221085 281311 221113
rect 281097 221023 281125 221051
rect 281159 221023 281187 221051
rect 281221 221023 281249 221051
rect 281283 221023 281311 221051
rect 281097 220961 281125 220989
rect 281159 220961 281187 220989
rect 281221 220961 281249 220989
rect 281283 220961 281311 220989
rect 281097 212147 281125 212175
rect 281159 212147 281187 212175
rect 281221 212147 281249 212175
rect 281283 212147 281311 212175
rect 281097 212085 281125 212113
rect 281159 212085 281187 212113
rect 281221 212085 281249 212113
rect 281283 212085 281311 212113
rect 281097 212023 281125 212051
rect 281159 212023 281187 212051
rect 281221 212023 281249 212051
rect 281283 212023 281311 212051
rect 281097 211961 281125 211989
rect 281159 211961 281187 211989
rect 281221 211961 281249 211989
rect 281283 211961 281311 211989
rect 281097 203147 281125 203175
rect 281159 203147 281187 203175
rect 281221 203147 281249 203175
rect 281283 203147 281311 203175
rect 281097 203085 281125 203113
rect 281159 203085 281187 203113
rect 281221 203085 281249 203113
rect 281283 203085 281311 203113
rect 281097 203023 281125 203051
rect 281159 203023 281187 203051
rect 281221 203023 281249 203051
rect 281283 203023 281311 203051
rect 281097 202961 281125 202989
rect 281159 202961 281187 202989
rect 281221 202961 281249 202989
rect 281283 202961 281311 202989
rect 281097 194147 281125 194175
rect 281159 194147 281187 194175
rect 281221 194147 281249 194175
rect 281283 194147 281311 194175
rect 281097 194085 281125 194113
rect 281159 194085 281187 194113
rect 281221 194085 281249 194113
rect 281283 194085 281311 194113
rect 281097 194023 281125 194051
rect 281159 194023 281187 194051
rect 281221 194023 281249 194051
rect 281283 194023 281311 194051
rect 281097 193961 281125 193989
rect 281159 193961 281187 193989
rect 281221 193961 281249 193989
rect 281283 193961 281311 193989
rect 281097 185147 281125 185175
rect 281159 185147 281187 185175
rect 281221 185147 281249 185175
rect 281283 185147 281311 185175
rect 281097 185085 281125 185113
rect 281159 185085 281187 185113
rect 281221 185085 281249 185113
rect 281283 185085 281311 185113
rect 281097 185023 281125 185051
rect 281159 185023 281187 185051
rect 281221 185023 281249 185051
rect 281283 185023 281311 185051
rect 281097 184961 281125 184989
rect 281159 184961 281187 184989
rect 281221 184961 281249 184989
rect 281283 184961 281311 184989
rect 281097 176147 281125 176175
rect 281159 176147 281187 176175
rect 281221 176147 281249 176175
rect 281283 176147 281311 176175
rect 281097 176085 281125 176113
rect 281159 176085 281187 176113
rect 281221 176085 281249 176113
rect 281283 176085 281311 176113
rect 281097 176023 281125 176051
rect 281159 176023 281187 176051
rect 281221 176023 281249 176051
rect 281283 176023 281311 176051
rect 281097 175961 281125 175989
rect 281159 175961 281187 175989
rect 281221 175961 281249 175989
rect 281283 175961 281311 175989
rect 281097 167147 281125 167175
rect 281159 167147 281187 167175
rect 281221 167147 281249 167175
rect 281283 167147 281311 167175
rect 281097 167085 281125 167113
rect 281159 167085 281187 167113
rect 281221 167085 281249 167113
rect 281283 167085 281311 167113
rect 281097 167023 281125 167051
rect 281159 167023 281187 167051
rect 281221 167023 281249 167051
rect 281283 167023 281311 167051
rect 281097 166961 281125 166989
rect 281159 166961 281187 166989
rect 281221 166961 281249 166989
rect 281283 166961 281311 166989
rect 281097 158147 281125 158175
rect 281159 158147 281187 158175
rect 281221 158147 281249 158175
rect 281283 158147 281311 158175
rect 281097 158085 281125 158113
rect 281159 158085 281187 158113
rect 281221 158085 281249 158113
rect 281283 158085 281311 158113
rect 281097 158023 281125 158051
rect 281159 158023 281187 158051
rect 281221 158023 281249 158051
rect 281283 158023 281311 158051
rect 281097 157961 281125 157989
rect 281159 157961 281187 157989
rect 281221 157961 281249 157989
rect 281283 157961 281311 157989
rect 294597 272147 294625 272175
rect 294659 272147 294687 272175
rect 294721 272147 294749 272175
rect 294783 272147 294811 272175
rect 294597 272085 294625 272113
rect 294659 272085 294687 272113
rect 294721 272085 294749 272113
rect 294783 272085 294811 272113
rect 294597 272023 294625 272051
rect 294659 272023 294687 272051
rect 294721 272023 294749 272051
rect 294783 272023 294811 272051
rect 294597 271961 294625 271989
rect 294659 271961 294687 271989
rect 294721 271961 294749 271989
rect 294783 271961 294811 271989
rect 281097 149147 281125 149175
rect 281159 149147 281187 149175
rect 281221 149147 281249 149175
rect 281283 149147 281311 149175
rect 281097 149085 281125 149113
rect 281159 149085 281187 149113
rect 281221 149085 281249 149113
rect 281283 149085 281311 149113
rect 281097 149023 281125 149051
rect 281159 149023 281187 149051
rect 281221 149023 281249 149051
rect 281283 149023 281311 149051
rect 281097 148961 281125 148989
rect 281159 148961 281187 148989
rect 281221 148961 281249 148989
rect 281283 148961 281311 148989
rect 281097 140147 281125 140175
rect 281159 140147 281187 140175
rect 281221 140147 281249 140175
rect 281283 140147 281311 140175
rect 281097 140085 281125 140113
rect 281159 140085 281187 140113
rect 281221 140085 281249 140113
rect 281283 140085 281311 140113
rect 281097 140023 281125 140051
rect 281159 140023 281187 140051
rect 281221 140023 281249 140051
rect 281283 140023 281311 140051
rect 281097 139961 281125 139989
rect 281159 139961 281187 139989
rect 281221 139961 281249 139989
rect 281283 139961 281311 139989
rect 281097 131147 281125 131175
rect 281159 131147 281187 131175
rect 281221 131147 281249 131175
rect 281283 131147 281311 131175
rect 281097 131085 281125 131113
rect 281159 131085 281187 131113
rect 281221 131085 281249 131113
rect 281283 131085 281311 131113
rect 281097 131023 281125 131051
rect 281159 131023 281187 131051
rect 281221 131023 281249 131051
rect 281283 131023 281311 131051
rect 281097 130961 281125 130989
rect 281159 130961 281187 130989
rect 281221 130961 281249 130989
rect 281283 130961 281311 130989
rect 281097 122147 281125 122175
rect 281159 122147 281187 122175
rect 281221 122147 281249 122175
rect 281283 122147 281311 122175
rect 281097 122085 281125 122113
rect 281159 122085 281187 122113
rect 281221 122085 281249 122113
rect 281283 122085 281311 122113
rect 281097 122023 281125 122051
rect 281159 122023 281187 122051
rect 281221 122023 281249 122051
rect 281283 122023 281311 122051
rect 281097 121961 281125 121989
rect 281159 121961 281187 121989
rect 281221 121961 281249 121989
rect 281283 121961 281311 121989
rect 281097 113147 281125 113175
rect 281159 113147 281187 113175
rect 281221 113147 281249 113175
rect 281283 113147 281311 113175
rect 281097 113085 281125 113113
rect 281159 113085 281187 113113
rect 281221 113085 281249 113113
rect 281283 113085 281311 113113
rect 281097 113023 281125 113051
rect 281159 113023 281187 113051
rect 281221 113023 281249 113051
rect 281283 113023 281311 113051
rect 281097 112961 281125 112989
rect 281159 112961 281187 112989
rect 281221 112961 281249 112989
rect 281283 112961 281311 112989
rect 294597 263147 294625 263175
rect 294659 263147 294687 263175
rect 294721 263147 294749 263175
rect 294783 263147 294811 263175
rect 294597 263085 294625 263113
rect 294659 263085 294687 263113
rect 294721 263085 294749 263113
rect 294783 263085 294811 263113
rect 294597 263023 294625 263051
rect 294659 263023 294687 263051
rect 294721 263023 294749 263051
rect 294783 263023 294811 263051
rect 294597 262961 294625 262989
rect 294659 262961 294687 262989
rect 294721 262961 294749 262989
rect 294783 262961 294811 262989
rect 294597 254147 294625 254175
rect 294659 254147 294687 254175
rect 294721 254147 294749 254175
rect 294783 254147 294811 254175
rect 294597 254085 294625 254113
rect 294659 254085 294687 254113
rect 294721 254085 294749 254113
rect 294783 254085 294811 254113
rect 294597 254023 294625 254051
rect 294659 254023 294687 254051
rect 294721 254023 294749 254051
rect 294783 254023 294811 254051
rect 294597 253961 294625 253989
rect 294659 253961 294687 253989
rect 294721 253961 294749 253989
rect 294783 253961 294811 253989
rect 281097 104147 281125 104175
rect 281159 104147 281187 104175
rect 281221 104147 281249 104175
rect 281283 104147 281311 104175
rect 281097 104085 281125 104113
rect 281159 104085 281187 104113
rect 281221 104085 281249 104113
rect 281283 104085 281311 104113
rect 281097 104023 281125 104051
rect 281159 104023 281187 104051
rect 281221 104023 281249 104051
rect 281283 104023 281311 104051
rect 281097 103961 281125 103989
rect 281159 103961 281187 103989
rect 281221 103961 281249 103989
rect 281283 103961 281311 103989
rect 281097 95147 281125 95175
rect 281159 95147 281187 95175
rect 281221 95147 281249 95175
rect 281283 95147 281311 95175
rect 281097 95085 281125 95113
rect 281159 95085 281187 95113
rect 281221 95085 281249 95113
rect 281283 95085 281311 95113
rect 281097 95023 281125 95051
rect 281159 95023 281187 95051
rect 281221 95023 281249 95051
rect 281283 95023 281311 95051
rect 281097 94961 281125 94989
rect 281159 94961 281187 94989
rect 281221 94961 281249 94989
rect 281283 94961 281311 94989
rect 281097 86147 281125 86175
rect 281159 86147 281187 86175
rect 281221 86147 281249 86175
rect 281283 86147 281311 86175
rect 281097 86085 281125 86113
rect 281159 86085 281187 86113
rect 281221 86085 281249 86113
rect 281283 86085 281311 86113
rect 281097 86023 281125 86051
rect 281159 86023 281187 86051
rect 281221 86023 281249 86051
rect 281283 86023 281311 86051
rect 281097 85961 281125 85989
rect 281159 85961 281187 85989
rect 281221 85961 281249 85989
rect 281283 85961 281311 85989
rect 281097 77147 281125 77175
rect 281159 77147 281187 77175
rect 281221 77147 281249 77175
rect 281283 77147 281311 77175
rect 281097 77085 281125 77113
rect 281159 77085 281187 77113
rect 281221 77085 281249 77113
rect 281283 77085 281311 77113
rect 281097 77023 281125 77051
rect 281159 77023 281187 77051
rect 281221 77023 281249 77051
rect 281283 77023 281311 77051
rect 281097 76961 281125 76989
rect 281159 76961 281187 76989
rect 281221 76961 281249 76989
rect 281283 76961 281311 76989
rect 281097 68147 281125 68175
rect 281159 68147 281187 68175
rect 281221 68147 281249 68175
rect 281283 68147 281311 68175
rect 281097 68085 281125 68113
rect 281159 68085 281187 68113
rect 281221 68085 281249 68113
rect 281283 68085 281311 68113
rect 281097 68023 281125 68051
rect 281159 68023 281187 68051
rect 281221 68023 281249 68051
rect 281283 68023 281311 68051
rect 281097 67961 281125 67989
rect 281159 67961 281187 67989
rect 281221 67961 281249 67989
rect 281283 67961 281311 67989
rect 281097 59147 281125 59175
rect 281159 59147 281187 59175
rect 281221 59147 281249 59175
rect 281283 59147 281311 59175
rect 281097 59085 281125 59113
rect 281159 59085 281187 59113
rect 281221 59085 281249 59113
rect 281283 59085 281311 59113
rect 281097 59023 281125 59051
rect 281159 59023 281187 59051
rect 281221 59023 281249 59051
rect 281283 59023 281311 59051
rect 281097 58961 281125 58989
rect 281159 58961 281187 58989
rect 281221 58961 281249 58989
rect 281283 58961 281311 58989
rect 281097 50147 281125 50175
rect 281159 50147 281187 50175
rect 281221 50147 281249 50175
rect 281283 50147 281311 50175
rect 281097 50085 281125 50113
rect 281159 50085 281187 50113
rect 281221 50085 281249 50113
rect 281283 50085 281311 50113
rect 281097 50023 281125 50051
rect 281159 50023 281187 50051
rect 281221 50023 281249 50051
rect 281283 50023 281311 50051
rect 281097 49961 281125 49989
rect 281159 49961 281187 49989
rect 281221 49961 281249 49989
rect 281283 49961 281311 49989
rect 281097 41147 281125 41175
rect 281159 41147 281187 41175
rect 281221 41147 281249 41175
rect 281283 41147 281311 41175
rect 281097 41085 281125 41113
rect 281159 41085 281187 41113
rect 281221 41085 281249 41113
rect 281283 41085 281311 41113
rect 281097 41023 281125 41051
rect 281159 41023 281187 41051
rect 281221 41023 281249 41051
rect 281283 41023 281311 41051
rect 281097 40961 281125 40989
rect 281159 40961 281187 40989
rect 281221 40961 281249 40989
rect 281283 40961 281311 40989
rect 281097 32147 281125 32175
rect 281159 32147 281187 32175
rect 281221 32147 281249 32175
rect 281283 32147 281311 32175
rect 281097 32085 281125 32113
rect 281159 32085 281187 32113
rect 281221 32085 281249 32113
rect 281283 32085 281311 32113
rect 281097 32023 281125 32051
rect 281159 32023 281187 32051
rect 281221 32023 281249 32051
rect 281283 32023 281311 32051
rect 281097 31961 281125 31989
rect 281159 31961 281187 31989
rect 281221 31961 281249 31989
rect 281283 31961 281311 31989
rect 281097 23147 281125 23175
rect 281159 23147 281187 23175
rect 281221 23147 281249 23175
rect 281283 23147 281311 23175
rect 281097 23085 281125 23113
rect 281159 23085 281187 23113
rect 281221 23085 281249 23113
rect 281283 23085 281311 23113
rect 281097 23023 281125 23051
rect 281159 23023 281187 23051
rect 281221 23023 281249 23051
rect 281283 23023 281311 23051
rect 281097 22961 281125 22989
rect 281159 22961 281187 22989
rect 281221 22961 281249 22989
rect 281283 22961 281311 22989
rect 281097 14147 281125 14175
rect 281159 14147 281187 14175
rect 281221 14147 281249 14175
rect 281283 14147 281311 14175
rect 281097 14085 281125 14113
rect 281159 14085 281187 14113
rect 281221 14085 281249 14113
rect 281283 14085 281311 14113
rect 281097 14023 281125 14051
rect 281159 14023 281187 14051
rect 281221 14023 281249 14051
rect 281283 14023 281311 14051
rect 281097 13961 281125 13989
rect 281159 13961 281187 13989
rect 281221 13961 281249 13989
rect 281283 13961 281311 13989
rect 281097 5147 281125 5175
rect 281159 5147 281187 5175
rect 281221 5147 281249 5175
rect 281283 5147 281311 5175
rect 281097 5085 281125 5113
rect 281159 5085 281187 5113
rect 281221 5085 281249 5113
rect 281283 5085 281311 5113
rect 281097 5023 281125 5051
rect 281159 5023 281187 5051
rect 281221 5023 281249 5051
rect 281283 5023 281311 5051
rect 281097 4961 281125 4989
rect 281159 4961 281187 4989
rect 281221 4961 281249 4989
rect 281283 4961 281311 4989
rect 294597 245147 294625 245175
rect 294659 245147 294687 245175
rect 294721 245147 294749 245175
rect 294783 245147 294811 245175
rect 294597 245085 294625 245113
rect 294659 245085 294687 245113
rect 294721 245085 294749 245113
rect 294783 245085 294811 245113
rect 294597 245023 294625 245051
rect 294659 245023 294687 245051
rect 294721 245023 294749 245051
rect 294783 245023 294811 245051
rect 294597 244961 294625 244989
rect 294659 244961 294687 244989
rect 294721 244961 294749 244989
rect 294783 244961 294811 244989
rect 294597 236147 294625 236175
rect 294659 236147 294687 236175
rect 294721 236147 294749 236175
rect 294783 236147 294811 236175
rect 294597 236085 294625 236113
rect 294659 236085 294687 236113
rect 294721 236085 294749 236113
rect 294783 236085 294811 236113
rect 294597 236023 294625 236051
rect 294659 236023 294687 236051
rect 294721 236023 294749 236051
rect 294783 236023 294811 236051
rect 294597 235961 294625 235989
rect 294659 235961 294687 235989
rect 294721 235961 294749 235989
rect 294783 235961 294811 235989
rect 294597 227147 294625 227175
rect 294659 227147 294687 227175
rect 294721 227147 294749 227175
rect 294783 227147 294811 227175
rect 294597 227085 294625 227113
rect 294659 227085 294687 227113
rect 294721 227085 294749 227113
rect 294783 227085 294811 227113
rect 294597 227023 294625 227051
rect 294659 227023 294687 227051
rect 294721 227023 294749 227051
rect 294783 227023 294811 227051
rect 294597 226961 294625 226989
rect 294659 226961 294687 226989
rect 294721 226961 294749 226989
rect 294783 226961 294811 226989
rect 294597 218147 294625 218175
rect 294659 218147 294687 218175
rect 294721 218147 294749 218175
rect 294783 218147 294811 218175
rect 294597 218085 294625 218113
rect 294659 218085 294687 218113
rect 294721 218085 294749 218113
rect 294783 218085 294811 218113
rect 294597 218023 294625 218051
rect 294659 218023 294687 218051
rect 294721 218023 294749 218051
rect 294783 218023 294811 218051
rect 294597 217961 294625 217989
rect 294659 217961 294687 217989
rect 294721 217961 294749 217989
rect 294783 217961 294811 217989
rect 294597 209147 294625 209175
rect 294659 209147 294687 209175
rect 294721 209147 294749 209175
rect 294783 209147 294811 209175
rect 294597 209085 294625 209113
rect 294659 209085 294687 209113
rect 294721 209085 294749 209113
rect 294783 209085 294811 209113
rect 294597 209023 294625 209051
rect 294659 209023 294687 209051
rect 294721 209023 294749 209051
rect 294783 209023 294811 209051
rect 294597 208961 294625 208989
rect 294659 208961 294687 208989
rect 294721 208961 294749 208989
rect 294783 208961 294811 208989
rect 294597 200147 294625 200175
rect 294659 200147 294687 200175
rect 294721 200147 294749 200175
rect 294783 200147 294811 200175
rect 294597 200085 294625 200113
rect 294659 200085 294687 200113
rect 294721 200085 294749 200113
rect 294783 200085 294811 200113
rect 294597 200023 294625 200051
rect 294659 200023 294687 200051
rect 294721 200023 294749 200051
rect 294783 200023 294811 200051
rect 294597 199961 294625 199989
rect 294659 199961 294687 199989
rect 294721 199961 294749 199989
rect 294783 199961 294811 199989
rect 294597 191147 294625 191175
rect 294659 191147 294687 191175
rect 294721 191147 294749 191175
rect 294783 191147 294811 191175
rect 294597 191085 294625 191113
rect 294659 191085 294687 191113
rect 294721 191085 294749 191113
rect 294783 191085 294811 191113
rect 294597 191023 294625 191051
rect 294659 191023 294687 191051
rect 294721 191023 294749 191051
rect 294783 191023 294811 191051
rect 294597 190961 294625 190989
rect 294659 190961 294687 190989
rect 294721 190961 294749 190989
rect 294783 190961 294811 190989
rect 294597 182147 294625 182175
rect 294659 182147 294687 182175
rect 294721 182147 294749 182175
rect 294783 182147 294811 182175
rect 294597 182085 294625 182113
rect 294659 182085 294687 182113
rect 294721 182085 294749 182113
rect 294783 182085 294811 182113
rect 294597 182023 294625 182051
rect 294659 182023 294687 182051
rect 294721 182023 294749 182051
rect 294783 182023 294811 182051
rect 294597 181961 294625 181989
rect 294659 181961 294687 181989
rect 294721 181961 294749 181989
rect 294783 181961 294811 181989
rect 294597 173147 294625 173175
rect 294659 173147 294687 173175
rect 294721 173147 294749 173175
rect 294783 173147 294811 173175
rect 294597 173085 294625 173113
rect 294659 173085 294687 173113
rect 294721 173085 294749 173113
rect 294783 173085 294811 173113
rect 294597 173023 294625 173051
rect 294659 173023 294687 173051
rect 294721 173023 294749 173051
rect 294783 173023 294811 173051
rect 294597 172961 294625 172989
rect 294659 172961 294687 172989
rect 294721 172961 294749 172989
rect 294783 172961 294811 172989
rect 294597 164147 294625 164175
rect 294659 164147 294687 164175
rect 294721 164147 294749 164175
rect 294783 164147 294811 164175
rect 294597 164085 294625 164113
rect 294659 164085 294687 164113
rect 294721 164085 294749 164113
rect 294783 164085 294811 164113
rect 294597 164023 294625 164051
rect 294659 164023 294687 164051
rect 294721 164023 294749 164051
rect 294783 164023 294811 164051
rect 294597 163961 294625 163989
rect 294659 163961 294687 163989
rect 294721 163961 294749 163989
rect 294783 163961 294811 163989
rect 294597 155147 294625 155175
rect 294659 155147 294687 155175
rect 294721 155147 294749 155175
rect 294783 155147 294811 155175
rect 294597 155085 294625 155113
rect 294659 155085 294687 155113
rect 294721 155085 294749 155113
rect 294783 155085 294811 155113
rect 294597 155023 294625 155051
rect 294659 155023 294687 155051
rect 294721 155023 294749 155051
rect 294783 155023 294811 155051
rect 294597 154961 294625 154989
rect 294659 154961 294687 154989
rect 294721 154961 294749 154989
rect 294783 154961 294811 154989
rect 294597 146147 294625 146175
rect 294659 146147 294687 146175
rect 294721 146147 294749 146175
rect 294783 146147 294811 146175
rect 294597 146085 294625 146113
rect 294659 146085 294687 146113
rect 294721 146085 294749 146113
rect 294783 146085 294811 146113
rect 294597 146023 294625 146051
rect 294659 146023 294687 146051
rect 294721 146023 294749 146051
rect 294783 146023 294811 146051
rect 294597 145961 294625 145989
rect 294659 145961 294687 145989
rect 294721 145961 294749 145989
rect 294783 145961 294811 145989
rect 294597 137147 294625 137175
rect 294659 137147 294687 137175
rect 294721 137147 294749 137175
rect 294783 137147 294811 137175
rect 294597 137085 294625 137113
rect 294659 137085 294687 137113
rect 294721 137085 294749 137113
rect 294783 137085 294811 137113
rect 294597 137023 294625 137051
rect 294659 137023 294687 137051
rect 294721 137023 294749 137051
rect 294783 137023 294811 137051
rect 294597 136961 294625 136989
rect 294659 136961 294687 136989
rect 294721 136961 294749 136989
rect 294783 136961 294811 136989
rect 294597 128147 294625 128175
rect 294659 128147 294687 128175
rect 294721 128147 294749 128175
rect 294783 128147 294811 128175
rect 294597 128085 294625 128113
rect 294659 128085 294687 128113
rect 294721 128085 294749 128113
rect 294783 128085 294811 128113
rect 294597 128023 294625 128051
rect 294659 128023 294687 128051
rect 294721 128023 294749 128051
rect 294783 128023 294811 128051
rect 294597 127961 294625 127989
rect 294659 127961 294687 127989
rect 294721 127961 294749 127989
rect 294783 127961 294811 127989
rect 294597 119147 294625 119175
rect 294659 119147 294687 119175
rect 294721 119147 294749 119175
rect 294783 119147 294811 119175
rect 294597 119085 294625 119113
rect 294659 119085 294687 119113
rect 294721 119085 294749 119113
rect 294783 119085 294811 119113
rect 294597 119023 294625 119051
rect 294659 119023 294687 119051
rect 294721 119023 294749 119051
rect 294783 119023 294811 119051
rect 294597 118961 294625 118989
rect 294659 118961 294687 118989
rect 294721 118961 294749 118989
rect 294783 118961 294811 118989
rect 294597 110147 294625 110175
rect 294659 110147 294687 110175
rect 294721 110147 294749 110175
rect 294783 110147 294811 110175
rect 294597 110085 294625 110113
rect 294659 110085 294687 110113
rect 294721 110085 294749 110113
rect 294783 110085 294811 110113
rect 294597 110023 294625 110051
rect 294659 110023 294687 110051
rect 294721 110023 294749 110051
rect 294783 110023 294811 110051
rect 294597 109961 294625 109989
rect 294659 109961 294687 109989
rect 294721 109961 294749 109989
rect 294783 109961 294811 109989
rect 294597 101147 294625 101175
rect 294659 101147 294687 101175
rect 294721 101147 294749 101175
rect 294783 101147 294811 101175
rect 294597 101085 294625 101113
rect 294659 101085 294687 101113
rect 294721 101085 294749 101113
rect 294783 101085 294811 101113
rect 294597 101023 294625 101051
rect 294659 101023 294687 101051
rect 294721 101023 294749 101051
rect 294783 101023 294811 101051
rect 294597 100961 294625 100989
rect 294659 100961 294687 100989
rect 294721 100961 294749 100989
rect 294783 100961 294811 100989
rect 294597 92147 294625 92175
rect 294659 92147 294687 92175
rect 294721 92147 294749 92175
rect 294783 92147 294811 92175
rect 294597 92085 294625 92113
rect 294659 92085 294687 92113
rect 294721 92085 294749 92113
rect 294783 92085 294811 92113
rect 294597 92023 294625 92051
rect 294659 92023 294687 92051
rect 294721 92023 294749 92051
rect 294783 92023 294811 92051
rect 294597 91961 294625 91989
rect 294659 91961 294687 91989
rect 294721 91961 294749 91989
rect 294783 91961 294811 91989
rect 294597 83147 294625 83175
rect 294659 83147 294687 83175
rect 294721 83147 294749 83175
rect 294783 83147 294811 83175
rect 294597 83085 294625 83113
rect 294659 83085 294687 83113
rect 294721 83085 294749 83113
rect 294783 83085 294811 83113
rect 294597 83023 294625 83051
rect 294659 83023 294687 83051
rect 294721 83023 294749 83051
rect 294783 83023 294811 83051
rect 294597 82961 294625 82989
rect 294659 82961 294687 82989
rect 294721 82961 294749 82989
rect 294783 82961 294811 82989
rect 294597 74147 294625 74175
rect 294659 74147 294687 74175
rect 294721 74147 294749 74175
rect 294783 74147 294811 74175
rect 294597 74085 294625 74113
rect 294659 74085 294687 74113
rect 294721 74085 294749 74113
rect 294783 74085 294811 74113
rect 294597 74023 294625 74051
rect 294659 74023 294687 74051
rect 294721 74023 294749 74051
rect 294783 74023 294811 74051
rect 294597 73961 294625 73989
rect 294659 73961 294687 73989
rect 294721 73961 294749 73989
rect 294783 73961 294811 73989
rect 294597 65147 294625 65175
rect 294659 65147 294687 65175
rect 294721 65147 294749 65175
rect 294783 65147 294811 65175
rect 294597 65085 294625 65113
rect 294659 65085 294687 65113
rect 294721 65085 294749 65113
rect 294783 65085 294811 65113
rect 294597 65023 294625 65051
rect 294659 65023 294687 65051
rect 294721 65023 294749 65051
rect 294783 65023 294811 65051
rect 294597 64961 294625 64989
rect 294659 64961 294687 64989
rect 294721 64961 294749 64989
rect 294783 64961 294811 64989
rect 294597 56147 294625 56175
rect 294659 56147 294687 56175
rect 294721 56147 294749 56175
rect 294783 56147 294811 56175
rect 294597 56085 294625 56113
rect 294659 56085 294687 56113
rect 294721 56085 294749 56113
rect 294783 56085 294811 56113
rect 294597 56023 294625 56051
rect 294659 56023 294687 56051
rect 294721 56023 294749 56051
rect 294783 56023 294811 56051
rect 294597 55961 294625 55989
rect 294659 55961 294687 55989
rect 294721 55961 294749 55989
rect 294783 55961 294811 55989
rect 294597 47147 294625 47175
rect 294659 47147 294687 47175
rect 294721 47147 294749 47175
rect 294783 47147 294811 47175
rect 294597 47085 294625 47113
rect 294659 47085 294687 47113
rect 294721 47085 294749 47113
rect 294783 47085 294811 47113
rect 294597 47023 294625 47051
rect 294659 47023 294687 47051
rect 294721 47023 294749 47051
rect 294783 47023 294811 47051
rect 294597 46961 294625 46989
rect 294659 46961 294687 46989
rect 294721 46961 294749 46989
rect 294783 46961 294811 46989
rect 294597 38147 294625 38175
rect 294659 38147 294687 38175
rect 294721 38147 294749 38175
rect 294783 38147 294811 38175
rect 294597 38085 294625 38113
rect 294659 38085 294687 38113
rect 294721 38085 294749 38113
rect 294783 38085 294811 38113
rect 294597 38023 294625 38051
rect 294659 38023 294687 38051
rect 294721 38023 294749 38051
rect 294783 38023 294811 38051
rect 294597 37961 294625 37989
rect 294659 37961 294687 37989
rect 294721 37961 294749 37989
rect 294783 37961 294811 37989
rect 294597 29147 294625 29175
rect 294659 29147 294687 29175
rect 294721 29147 294749 29175
rect 294783 29147 294811 29175
rect 294597 29085 294625 29113
rect 294659 29085 294687 29113
rect 294721 29085 294749 29113
rect 294783 29085 294811 29113
rect 294597 29023 294625 29051
rect 294659 29023 294687 29051
rect 294721 29023 294749 29051
rect 294783 29023 294811 29051
rect 294597 28961 294625 28989
rect 294659 28961 294687 28989
rect 294721 28961 294749 28989
rect 294783 28961 294811 28989
rect 294597 20147 294625 20175
rect 294659 20147 294687 20175
rect 294721 20147 294749 20175
rect 294783 20147 294811 20175
rect 294597 20085 294625 20113
rect 294659 20085 294687 20113
rect 294721 20085 294749 20113
rect 294783 20085 294811 20113
rect 294597 20023 294625 20051
rect 294659 20023 294687 20051
rect 294721 20023 294749 20051
rect 294783 20023 294811 20051
rect 294597 19961 294625 19989
rect 294659 19961 294687 19989
rect 294721 19961 294749 19989
rect 294783 19961 294811 19989
rect 294597 11147 294625 11175
rect 294659 11147 294687 11175
rect 294721 11147 294749 11175
rect 294783 11147 294811 11175
rect 294597 11085 294625 11113
rect 294659 11085 294687 11113
rect 294721 11085 294749 11113
rect 294783 11085 294811 11113
rect 294597 11023 294625 11051
rect 294659 11023 294687 11051
rect 294721 11023 294749 11051
rect 294783 11023 294811 11051
rect 294597 10961 294625 10989
rect 294659 10961 294687 10989
rect 294721 10961 294749 10989
rect 294783 10961 294811 10989
rect 281097 -588 281125 -560
rect 281159 -588 281187 -560
rect 281221 -588 281249 -560
rect 281283 -588 281311 -560
rect 281097 -650 281125 -622
rect 281159 -650 281187 -622
rect 281221 -650 281249 -622
rect 281283 -650 281311 -622
rect 281097 -712 281125 -684
rect 281159 -712 281187 -684
rect 281221 -712 281249 -684
rect 281283 -712 281311 -684
rect 281097 -774 281125 -746
rect 281159 -774 281187 -746
rect 281221 -774 281249 -746
rect 281283 -774 281311 -746
rect 294597 2147 294625 2175
rect 294659 2147 294687 2175
rect 294721 2147 294749 2175
rect 294783 2147 294811 2175
rect 294597 2085 294625 2113
rect 294659 2085 294687 2113
rect 294721 2085 294749 2113
rect 294783 2085 294811 2113
rect 294597 2023 294625 2051
rect 294659 2023 294687 2051
rect 294721 2023 294749 2051
rect 294783 2023 294811 2051
rect 294597 1961 294625 1989
rect 294659 1961 294687 1989
rect 294721 1961 294749 1989
rect 294783 1961 294811 1989
rect 294597 -108 294625 -80
rect 294659 -108 294687 -80
rect 294721 -108 294749 -80
rect 294783 -108 294811 -80
rect 294597 -170 294625 -142
rect 294659 -170 294687 -142
rect 294721 -170 294749 -142
rect 294783 -170 294811 -142
rect 294597 -232 294625 -204
rect 294659 -232 294687 -204
rect 294721 -232 294749 -204
rect 294783 -232 294811 -204
rect 294597 -294 294625 -266
rect 294659 -294 294687 -266
rect 294721 -294 294749 -266
rect 294783 -294 294811 -266
rect 296457 299058 296485 299086
rect 296519 299058 296547 299086
rect 296581 299058 296609 299086
rect 296643 299058 296671 299086
rect 296457 298996 296485 299024
rect 296519 298996 296547 299024
rect 296581 298996 296609 299024
rect 296643 298996 296671 299024
rect 296457 298934 296485 298962
rect 296519 298934 296547 298962
rect 296581 298934 296609 298962
rect 296643 298934 296671 298962
rect 296457 298872 296485 298900
rect 296519 298872 296547 298900
rect 296581 298872 296609 298900
rect 296643 298872 296671 298900
rect 298728 299058 298756 299086
rect 298790 299058 298818 299086
rect 298852 299058 298880 299086
rect 298914 299058 298942 299086
rect 298728 298996 298756 299024
rect 298790 298996 298818 299024
rect 298852 298996 298880 299024
rect 298914 298996 298942 299024
rect 298728 298934 298756 298962
rect 298790 298934 298818 298962
rect 298852 298934 298880 298962
rect 298914 298934 298942 298962
rect 298728 298872 298756 298900
rect 298790 298872 298818 298900
rect 298852 298872 298880 298900
rect 298914 298872 298942 298900
rect 296457 293147 296485 293175
rect 296519 293147 296547 293175
rect 296581 293147 296609 293175
rect 296643 293147 296671 293175
rect 296457 293085 296485 293113
rect 296519 293085 296547 293113
rect 296581 293085 296609 293113
rect 296643 293085 296671 293113
rect 296457 293023 296485 293051
rect 296519 293023 296547 293051
rect 296581 293023 296609 293051
rect 296643 293023 296671 293051
rect 296457 292961 296485 292989
rect 296519 292961 296547 292989
rect 296581 292961 296609 292989
rect 296643 292961 296671 292989
rect 296457 284147 296485 284175
rect 296519 284147 296547 284175
rect 296581 284147 296609 284175
rect 296643 284147 296671 284175
rect 296457 284085 296485 284113
rect 296519 284085 296547 284113
rect 296581 284085 296609 284113
rect 296643 284085 296671 284113
rect 296457 284023 296485 284051
rect 296519 284023 296547 284051
rect 296581 284023 296609 284051
rect 296643 284023 296671 284051
rect 296457 283961 296485 283989
rect 296519 283961 296547 283989
rect 296581 283961 296609 283989
rect 296643 283961 296671 283989
rect 296457 275147 296485 275175
rect 296519 275147 296547 275175
rect 296581 275147 296609 275175
rect 296643 275147 296671 275175
rect 296457 275085 296485 275113
rect 296519 275085 296547 275113
rect 296581 275085 296609 275113
rect 296643 275085 296671 275113
rect 296457 275023 296485 275051
rect 296519 275023 296547 275051
rect 296581 275023 296609 275051
rect 296643 275023 296671 275051
rect 296457 274961 296485 274989
rect 296519 274961 296547 274989
rect 296581 274961 296609 274989
rect 296643 274961 296671 274989
rect 296457 266147 296485 266175
rect 296519 266147 296547 266175
rect 296581 266147 296609 266175
rect 296643 266147 296671 266175
rect 296457 266085 296485 266113
rect 296519 266085 296547 266113
rect 296581 266085 296609 266113
rect 296643 266085 296671 266113
rect 296457 266023 296485 266051
rect 296519 266023 296547 266051
rect 296581 266023 296609 266051
rect 296643 266023 296671 266051
rect 296457 265961 296485 265989
rect 296519 265961 296547 265989
rect 296581 265961 296609 265989
rect 296643 265961 296671 265989
rect 296457 257147 296485 257175
rect 296519 257147 296547 257175
rect 296581 257147 296609 257175
rect 296643 257147 296671 257175
rect 296457 257085 296485 257113
rect 296519 257085 296547 257113
rect 296581 257085 296609 257113
rect 296643 257085 296671 257113
rect 296457 257023 296485 257051
rect 296519 257023 296547 257051
rect 296581 257023 296609 257051
rect 296643 257023 296671 257051
rect 296457 256961 296485 256989
rect 296519 256961 296547 256989
rect 296581 256961 296609 256989
rect 296643 256961 296671 256989
rect 296457 248147 296485 248175
rect 296519 248147 296547 248175
rect 296581 248147 296609 248175
rect 296643 248147 296671 248175
rect 296457 248085 296485 248113
rect 296519 248085 296547 248113
rect 296581 248085 296609 248113
rect 296643 248085 296671 248113
rect 296457 248023 296485 248051
rect 296519 248023 296547 248051
rect 296581 248023 296609 248051
rect 296643 248023 296671 248051
rect 296457 247961 296485 247989
rect 296519 247961 296547 247989
rect 296581 247961 296609 247989
rect 296643 247961 296671 247989
rect 296457 239147 296485 239175
rect 296519 239147 296547 239175
rect 296581 239147 296609 239175
rect 296643 239147 296671 239175
rect 296457 239085 296485 239113
rect 296519 239085 296547 239113
rect 296581 239085 296609 239113
rect 296643 239085 296671 239113
rect 296457 239023 296485 239051
rect 296519 239023 296547 239051
rect 296581 239023 296609 239051
rect 296643 239023 296671 239051
rect 296457 238961 296485 238989
rect 296519 238961 296547 238989
rect 296581 238961 296609 238989
rect 296643 238961 296671 238989
rect 296457 230147 296485 230175
rect 296519 230147 296547 230175
rect 296581 230147 296609 230175
rect 296643 230147 296671 230175
rect 296457 230085 296485 230113
rect 296519 230085 296547 230113
rect 296581 230085 296609 230113
rect 296643 230085 296671 230113
rect 296457 230023 296485 230051
rect 296519 230023 296547 230051
rect 296581 230023 296609 230051
rect 296643 230023 296671 230051
rect 296457 229961 296485 229989
rect 296519 229961 296547 229989
rect 296581 229961 296609 229989
rect 296643 229961 296671 229989
rect 296457 221147 296485 221175
rect 296519 221147 296547 221175
rect 296581 221147 296609 221175
rect 296643 221147 296671 221175
rect 296457 221085 296485 221113
rect 296519 221085 296547 221113
rect 296581 221085 296609 221113
rect 296643 221085 296671 221113
rect 296457 221023 296485 221051
rect 296519 221023 296547 221051
rect 296581 221023 296609 221051
rect 296643 221023 296671 221051
rect 296457 220961 296485 220989
rect 296519 220961 296547 220989
rect 296581 220961 296609 220989
rect 296643 220961 296671 220989
rect 296457 212147 296485 212175
rect 296519 212147 296547 212175
rect 296581 212147 296609 212175
rect 296643 212147 296671 212175
rect 296457 212085 296485 212113
rect 296519 212085 296547 212113
rect 296581 212085 296609 212113
rect 296643 212085 296671 212113
rect 296457 212023 296485 212051
rect 296519 212023 296547 212051
rect 296581 212023 296609 212051
rect 296643 212023 296671 212051
rect 296457 211961 296485 211989
rect 296519 211961 296547 211989
rect 296581 211961 296609 211989
rect 296643 211961 296671 211989
rect 296457 203147 296485 203175
rect 296519 203147 296547 203175
rect 296581 203147 296609 203175
rect 296643 203147 296671 203175
rect 296457 203085 296485 203113
rect 296519 203085 296547 203113
rect 296581 203085 296609 203113
rect 296643 203085 296671 203113
rect 296457 203023 296485 203051
rect 296519 203023 296547 203051
rect 296581 203023 296609 203051
rect 296643 203023 296671 203051
rect 296457 202961 296485 202989
rect 296519 202961 296547 202989
rect 296581 202961 296609 202989
rect 296643 202961 296671 202989
rect 296457 194147 296485 194175
rect 296519 194147 296547 194175
rect 296581 194147 296609 194175
rect 296643 194147 296671 194175
rect 296457 194085 296485 194113
rect 296519 194085 296547 194113
rect 296581 194085 296609 194113
rect 296643 194085 296671 194113
rect 296457 194023 296485 194051
rect 296519 194023 296547 194051
rect 296581 194023 296609 194051
rect 296643 194023 296671 194051
rect 296457 193961 296485 193989
rect 296519 193961 296547 193989
rect 296581 193961 296609 193989
rect 296643 193961 296671 193989
rect 296457 185147 296485 185175
rect 296519 185147 296547 185175
rect 296581 185147 296609 185175
rect 296643 185147 296671 185175
rect 296457 185085 296485 185113
rect 296519 185085 296547 185113
rect 296581 185085 296609 185113
rect 296643 185085 296671 185113
rect 296457 185023 296485 185051
rect 296519 185023 296547 185051
rect 296581 185023 296609 185051
rect 296643 185023 296671 185051
rect 296457 184961 296485 184989
rect 296519 184961 296547 184989
rect 296581 184961 296609 184989
rect 296643 184961 296671 184989
rect 296457 176147 296485 176175
rect 296519 176147 296547 176175
rect 296581 176147 296609 176175
rect 296643 176147 296671 176175
rect 296457 176085 296485 176113
rect 296519 176085 296547 176113
rect 296581 176085 296609 176113
rect 296643 176085 296671 176113
rect 296457 176023 296485 176051
rect 296519 176023 296547 176051
rect 296581 176023 296609 176051
rect 296643 176023 296671 176051
rect 296457 175961 296485 175989
rect 296519 175961 296547 175989
rect 296581 175961 296609 175989
rect 296643 175961 296671 175989
rect 296457 167147 296485 167175
rect 296519 167147 296547 167175
rect 296581 167147 296609 167175
rect 296643 167147 296671 167175
rect 296457 167085 296485 167113
rect 296519 167085 296547 167113
rect 296581 167085 296609 167113
rect 296643 167085 296671 167113
rect 296457 167023 296485 167051
rect 296519 167023 296547 167051
rect 296581 167023 296609 167051
rect 296643 167023 296671 167051
rect 296457 166961 296485 166989
rect 296519 166961 296547 166989
rect 296581 166961 296609 166989
rect 296643 166961 296671 166989
rect 296457 158147 296485 158175
rect 296519 158147 296547 158175
rect 296581 158147 296609 158175
rect 296643 158147 296671 158175
rect 296457 158085 296485 158113
rect 296519 158085 296547 158113
rect 296581 158085 296609 158113
rect 296643 158085 296671 158113
rect 296457 158023 296485 158051
rect 296519 158023 296547 158051
rect 296581 158023 296609 158051
rect 296643 158023 296671 158051
rect 296457 157961 296485 157989
rect 296519 157961 296547 157989
rect 296581 157961 296609 157989
rect 296643 157961 296671 157989
rect 296457 149147 296485 149175
rect 296519 149147 296547 149175
rect 296581 149147 296609 149175
rect 296643 149147 296671 149175
rect 296457 149085 296485 149113
rect 296519 149085 296547 149113
rect 296581 149085 296609 149113
rect 296643 149085 296671 149113
rect 296457 149023 296485 149051
rect 296519 149023 296547 149051
rect 296581 149023 296609 149051
rect 296643 149023 296671 149051
rect 296457 148961 296485 148989
rect 296519 148961 296547 148989
rect 296581 148961 296609 148989
rect 296643 148961 296671 148989
rect 296457 140147 296485 140175
rect 296519 140147 296547 140175
rect 296581 140147 296609 140175
rect 296643 140147 296671 140175
rect 296457 140085 296485 140113
rect 296519 140085 296547 140113
rect 296581 140085 296609 140113
rect 296643 140085 296671 140113
rect 296457 140023 296485 140051
rect 296519 140023 296547 140051
rect 296581 140023 296609 140051
rect 296643 140023 296671 140051
rect 296457 139961 296485 139989
rect 296519 139961 296547 139989
rect 296581 139961 296609 139989
rect 296643 139961 296671 139989
rect 296457 131147 296485 131175
rect 296519 131147 296547 131175
rect 296581 131147 296609 131175
rect 296643 131147 296671 131175
rect 296457 131085 296485 131113
rect 296519 131085 296547 131113
rect 296581 131085 296609 131113
rect 296643 131085 296671 131113
rect 296457 131023 296485 131051
rect 296519 131023 296547 131051
rect 296581 131023 296609 131051
rect 296643 131023 296671 131051
rect 296457 130961 296485 130989
rect 296519 130961 296547 130989
rect 296581 130961 296609 130989
rect 296643 130961 296671 130989
rect 296457 122147 296485 122175
rect 296519 122147 296547 122175
rect 296581 122147 296609 122175
rect 296643 122147 296671 122175
rect 296457 122085 296485 122113
rect 296519 122085 296547 122113
rect 296581 122085 296609 122113
rect 296643 122085 296671 122113
rect 296457 122023 296485 122051
rect 296519 122023 296547 122051
rect 296581 122023 296609 122051
rect 296643 122023 296671 122051
rect 296457 121961 296485 121989
rect 296519 121961 296547 121989
rect 296581 121961 296609 121989
rect 296643 121961 296671 121989
rect 296457 113147 296485 113175
rect 296519 113147 296547 113175
rect 296581 113147 296609 113175
rect 296643 113147 296671 113175
rect 296457 113085 296485 113113
rect 296519 113085 296547 113113
rect 296581 113085 296609 113113
rect 296643 113085 296671 113113
rect 296457 113023 296485 113051
rect 296519 113023 296547 113051
rect 296581 113023 296609 113051
rect 296643 113023 296671 113051
rect 296457 112961 296485 112989
rect 296519 112961 296547 112989
rect 296581 112961 296609 112989
rect 296643 112961 296671 112989
rect 296457 104147 296485 104175
rect 296519 104147 296547 104175
rect 296581 104147 296609 104175
rect 296643 104147 296671 104175
rect 296457 104085 296485 104113
rect 296519 104085 296547 104113
rect 296581 104085 296609 104113
rect 296643 104085 296671 104113
rect 296457 104023 296485 104051
rect 296519 104023 296547 104051
rect 296581 104023 296609 104051
rect 296643 104023 296671 104051
rect 296457 103961 296485 103989
rect 296519 103961 296547 103989
rect 296581 103961 296609 103989
rect 296643 103961 296671 103989
rect 296457 95147 296485 95175
rect 296519 95147 296547 95175
rect 296581 95147 296609 95175
rect 296643 95147 296671 95175
rect 296457 95085 296485 95113
rect 296519 95085 296547 95113
rect 296581 95085 296609 95113
rect 296643 95085 296671 95113
rect 296457 95023 296485 95051
rect 296519 95023 296547 95051
rect 296581 95023 296609 95051
rect 296643 95023 296671 95051
rect 296457 94961 296485 94989
rect 296519 94961 296547 94989
rect 296581 94961 296609 94989
rect 296643 94961 296671 94989
rect 296457 86147 296485 86175
rect 296519 86147 296547 86175
rect 296581 86147 296609 86175
rect 296643 86147 296671 86175
rect 296457 86085 296485 86113
rect 296519 86085 296547 86113
rect 296581 86085 296609 86113
rect 296643 86085 296671 86113
rect 296457 86023 296485 86051
rect 296519 86023 296547 86051
rect 296581 86023 296609 86051
rect 296643 86023 296671 86051
rect 296457 85961 296485 85989
rect 296519 85961 296547 85989
rect 296581 85961 296609 85989
rect 296643 85961 296671 85989
rect 296457 77147 296485 77175
rect 296519 77147 296547 77175
rect 296581 77147 296609 77175
rect 296643 77147 296671 77175
rect 296457 77085 296485 77113
rect 296519 77085 296547 77113
rect 296581 77085 296609 77113
rect 296643 77085 296671 77113
rect 296457 77023 296485 77051
rect 296519 77023 296547 77051
rect 296581 77023 296609 77051
rect 296643 77023 296671 77051
rect 296457 76961 296485 76989
rect 296519 76961 296547 76989
rect 296581 76961 296609 76989
rect 296643 76961 296671 76989
rect 296457 68147 296485 68175
rect 296519 68147 296547 68175
rect 296581 68147 296609 68175
rect 296643 68147 296671 68175
rect 296457 68085 296485 68113
rect 296519 68085 296547 68113
rect 296581 68085 296609 68113
rect 296643 68085 296671 68113
rect 296457 68023 296485 68051
rect 296519 68023 296547 68051
rect 296581 68023 296609 68051
rect 296643 68023 296671 68051
rect 296457 67961 296485 67989
rect 296519 67961 296547 67989
rect 296581 67961 296609 67989
rect 296643 67961 296671 67989
rect 296457 59147 296485 59175
rect 296519 59147 296547 59175
rect 296581 59147 296609 59175
rect 296643 59147 296671 59175
rect 296457 59085 296485 59113
rect 296519 59085 296547 59113
rect 296581 59085 296609 59113
rect 296643 59085 296671 59113
rect 296457 59023 296485 59051
rect 296519 59023 296547 59051
rect 296581 59023 296609 59051
rect 296643 59023 296671 59051
rect 296457 58961 296485 58989
rect 296519 58961 296547 58989
rect 296581 58961 296609 58989
rect 296643 58961 296671 58989
rect 296457 50147 296485 50175
rect 296519 50147 296547 50175
rect 296581 50147 296609 50175
rect 296643 50147 296671 50175
rect 296457 50085 296485 50113
rect 296519 50085 296547 50113
rect 296581 50085 296609 50113
rect 296643 50085 296671 50113
rect 296457 50023 296485 50051
rect 296519 50023 296547 50051
rect 296581 50023 296609 50051
rect 296643 50023 296671 50051
rect 296457 49961 296485 49989
rect 296519 49961 296547 49989
rect 296581 49961 296609 49989
rect 296643 49961 296671 49989
rect 296457 41147 296485 41175
rect 296519 41147 296547 41175
rect 296581 41147 296609 41175
rect 296643 41147 296671 41175
rect 296457 41085 296485 41113
rect 296519 41085 296547 41113
rect 296581 41085 296609 41113
rect 296643 41085 296671 41113
rect 296457 41023 296485 41051
rect 296519 41023 296547 41051
rect 296581 41023 296609 41051
rect 296643 41023 296671 41051
rect 296457 40961 296485 40989
rect 296519 40961 296547 40989
rect 296581 40961 296609 40989
rect 296643 40961 296671 40989
rect 296457 32147 296485 32175
rect 296519 32147 296547 32175
rect 296581 32147 296609 32175
rect 296643 32147 296671 32175
rect 296457 32085 296485 32113
rect 296519 32085 296547 32113
rect 296581 32085 296609 32113
rect 296643 32085 296671 32113
rect 296457 32023 296485 32051
rect 296519 32023 296547 32051
rect 296581 32023 296609 32051
rect 296643 32023 296671 32051
rect 296457 31961 296485 31989
rect 296519 31961 296547 31989
rect 296581 31961 296609 31989
rect 296643 31961 296671 31989
rect 296457 23147 296485 23175
rect 296519 23147 296547 23175
rect 296581 23147 296609 23175
rect 296643 23147 296671 23175
rect 296457 23085 296485 23113
rect 296519 23085 296547 23113
rect 296581 23085 296609 23113
rect 296643 23085 296671 23113
rect 296457 23023 296485 23051
rect 296519 23023 296547 23051
rect 296581 23023 296609 23051
rect 296643 23023 296671 23051
rect 296457 22961 296485 22989
rect 296519 22961 296547 22989
rect 296581 22961 296609 22989
rect 296643 22961 296671 22989
rect 296457 14147 296485 14175
rect 296519 14147 296547 14175
rect 296581 14147 296609 14175
rect 296643 14147 296671 14175
rect 296457 14085 296485 14113
rect 296519 14085 296547 14113
rect 296581 14085 296609 14113
rect 296643 14085 296671 14113
rect 296457 14023 296485 14051
rect 296519 14023 296547 14051
rect 296581 14023 296609 14051
rect 296643 14023 296671 14051
rect 296457 13961 296485 13989
rect 296519 13961 296547 13989
rect 296581 13961 296609 13989
rect 296643 13961 296671 13989
rect 296457 5147 296485 5175
rect 296519 5147 296547 5175
rect 296581 5147 296609 5175
rect 296643 5147 296671 5175
rect 296457 5085 296485 5113
rect 296519 5085 296547 5113
rect 296581 5085 296609 5113
rect 296643 5085 296671 5113
rect 296457 5023 296485 5051
rect 296519 5023 296547 5051
rect 296581 5023 296609 5051
rect 296643 5023 296671 5051
rect 296457 4961 296485 4989
rect 296519 4961 296547 4989
rect 296581 4961 296609 4989
rect 296643 4961 296671 4989
rect 298248 298578 298276 298606
rect 298310 298578 298338 298606
rect 298372 298578 298400 298606
rect 298434 298578 298462 298606
rect 298248 298516 298276 298544
rect 298310 298516 298338 298544
rect 298372 298516 298400 298544
rect 298434 298516 298462 298544
rect 298248 298454 298276 298482
rect 298310 298454 298338 298482
rect 298372 298454 298400 298482
rect 298434 298454 298462 298482
rect 298248 298392 298276 298420
rect 298310 298392 298338 298420
rect 298372 298392 298400 298420
rect 298434 298392 298462 298420
rect 298248 290147 298276 290175
rect 298310 290147 298338 290175
rect 298372 290147 298400 290175
rect 298434 290147 298462 290175
rect 298248 290085 298276 290113
rect 298310 290085 298338 290113
rect 298372 290085 298400 290113
rect 298434 290085 298462 290113
rect 298248 290023 298276 290051
rect 298310 290023 298338 290051
rect 298372 290023 298400 290051
rect 298434 290023 298462 290051
rect 298248 289961 298276 289989
rect 298310 289961 298338 289989
rect 298372 289961 298400 289989
rect 298434 289961 298462 289989
rect 298248 281147 298276 281175
rect 298310 281147 298338 281175
rect 298372 281147 298400 281175
rect 298434 281147 298462 281175
rect 298248 281085 298276 281113
rect 298310 281085 298338 281113
rect 298372 281085 298400 281113
rect 298434 281085 298462 281113
rect 298248 281023 298276 281051
rect 298310 281023 298338 281051
rect 298372 281023 298400 281051
rect 298434 281023 298462 281051
rect 298248 280961 298276 280989
rect 298310 280961 298338 280989
rect 298372 280961 298400 280989
rect 298434 280961 298462 280989
rect 298248 272147 298276 272175
rect 298310 272147 298338 272175
rect 298372 272147 298400 272175
rect 298434 272147 298462 272175
rect 298248 272085 298276 272113
rect 298310 272085 298338 272113
rect 298372 272085 298400 272113
rect 298434 272085 298462 272113
rect 298248 272023 298276 272051
rect 298310 272023 298338 272051
rect 298372 272023 298400 272051
rect 298434 272023 298462 272051
rect 298248 271961 298276 271989
rect 298310 271961 298338 271989
rect 298372 271961 298400 271989
rect 298434 271961 298462 271989
rect 298248 263147 298276 263175
rect 298310 263147 298338 263175
rect 298372 263147 298400 263175
rect 298434 263147 298462 263175
rect 298248 263085 298276 263113
rect 298310 263085 298338 263113
rect 298372 263085 298400 263113
rect 298434 263085 298462 263113
rect 298248 263023 298276 263051
rect 298310 263023 298338 263051
rect 298372 263023 298400 263051
rect 298434 263023 298462 263051
rect 298248 262961 298276 262989
rect 298310 262961 298338 262989
rect 298372 262961 298400 262989
rect 298434 262961 298462 262989
rect 298248 254147 298276 254175
rect 298310 254147 298338 254175
rect 298372 254147 298400 254175
rect 298434 254147 298462 254175
rect 298248 254085 298276 254113
rect 298310 254085 298338 254113
rect 298372 254085 298400 254113
rect 298434 254085 298462 254113
rect 298248 254023 298276 254051
rect 298310 254023 298338 254051
rect 298372 254023 298400 254051
rect 298434 254023 298462 254051
rect 298248 253961 298276 253989
rect 298310 253961 298338 253989
rect 298372 253961 298400 253989
rect 298434 253961 298462 253989
rect 298248 245147 298276 245175
rect 298310 245147 298338 245175
rect 298372 245147 298400 245175
rect 298434 245147 298462 245175
rect 298248 245085 298276 245113
rect 298310 245085 298338 245113
rect 298372 245085 298400 245113
rect 298434 245085 298462 245113
rect 298248 245023 298276 245051
rect 298310 245023 298338 245051
rect 298372 245023 298400 245051
rect 298434 245023 298462 245051
rect 298248 244961 298276 244989
rect 298310 244961 298338 244989
rect 298372 244961 298400 244989
rect 298434 244961 298462 244989
rect 298248 236147 298276 236175
rect 298310 236147 298338 236175
rect 298372 236147 298400 236175
rect 298434 236147 298462 236175
rect 298248 236085 298276 236113
rect 298310 236085 298338 236113
rect 298372 236085 298400 236113
rect 298434 236085 298462 236113
rect 298248 236023 298276 236051
rect 298310 236023 298338 236051
rect 298372 236023 298400 236051
rect 298434 236023 298462 236051
rect 298248 235961 298276 235989
rect 298310 235961 298338 235989
rect 298372 235961 298400 235989
rect 298434 235961 298462 235989
rect 298248 227147 298276 227175
rect 298310 227147 298338 227175
rect 298372 227147 298400 227175
rect 298434 227147 298462 227175
rect 298248 227085 298276 227113
rect 298310 227085 298338 227113
rect 298372 227085 298400 227113
rect 298434 227085 298462 227113
rect 298248 227023 298276 227051
rect 298310 227023 298338 227051
rect 298372 227023 298400 227051
rect 298434 227023 298462 227051
rect 298248 226961 298276 226989
rect 298310 226961 298338 226989
rect 298372 226961 298400 226989
rect 298434 226961 298462 226989
rect 298248 218147 298276 218175
rect 298310 218147 298338 218175
rect 298372 218147 298400 218175
rect 298434 218147 298462 218175
rect 298248 218085 298276 218113
rect 298310 218085 298338 218113
rect 298372 218085 298400 218113
rect 298434 218085 298462 218113
rect 298248 218023 298276 218051
rect 298310 218023 298338 218051
rect 298372 218023 298400 218051
rect 298434 218023 298462 218051
rect 298248 217961 298276 217989
rect 298310 217961 298338 217989
rect 298372 217961 298400 217989
rect 298434 217961 298462 217989
rect 298248 209147 298276 209175
rect 298310 209147 298338 209175
rect 298372 209147 298400 209175
rect 298434 209147 298462 209175
rect 298248 209085 298276 209113
rect 298310 209085 298338 209113
rect 298372 209085 298400 209113
rect 298434 209085 298462 209113
rect 298248 209023 298276 209051
rect 298310 209023 298338 209051
rect 298372 209023 298400 209051
rect 298434 209023 298462 209051
rect 298248 208961 298276 208989
rect 298310 208961 298338 208989
rect 298372 208961 298400 208989
rect 298434 208961 298462 208989
rect 298248 200147 298276 200175
rect 298310 200147 298338 200175
rect 298372 200147 298400 200175
rect 298434 200147 298462 200175
rect 298248 200085 298276 200113
rect 298310 200085 298338 200113
rect 298372 200085 298400 200113
rect 298434 200085 298462 200113
rect 298248 200023 298276 200051
rect 298310 200023 298338 200051
rect 298372 200023 298400 200051
rect 298434 200023 298462 200051
rect 298248 199961 298276 199989
rect 298310 199961 298338 199989
rect 298372 199961 298400 199989
rect 298434 199961 298462 199989
rect 298248 191147 298276 191175
rect 298310 191147 298338 191175
rect 298372 191147 298400 191175
rect 298434 191147 298462 191175
rect 298248 191085 298276 191113
rect 298310 191085 298338 191113
rect 298372 191085 298400 191113
rect 298434 191085 298462 191113
rect 298248 191023 298276 191051
rect 298310 191023 298338 191051
rect 298372 191023 298400 191051
rect 298434 191023 298462 191051
rect 298248 190961 298276 190989
rect 298310 190961 298338 190989
rect 298372 190961 298400 190989
rect 298434 190961 298462 190989
rect 298248 182147 298276 182175
rect 298310 182147 298338 182175
rect 298372 182147 298400 182175
rect 298434 182147 298462 182175
rect 298248 182085 298276 182113
rect 298310 182085 298338 182113
rect 298372 182085 298400 182113
rect 298434 182085 298462 182113
rect 298248 182023 298276 182051
rect 298310 182023 298338 182051
rect 298372 182023 298400 182051
rect 298434 182023 298462 182051
rect 298248 181961 298276 181989
rect 298310 181961 298338 181989
rect 298372 181961 298400 181989
rect 298434 181961 298462 181989
rect 298248 173147 298276 173175
rect 298310 173147 298338 173175
rect 298372 173147 298400 173175
rect 298434 173147 298462 173175
rect 298248 173085 298276 173113
rect 298310 173085 298338 173113
rect 298372 173085 298400 173113
rect 298434 173085 298462 173113
rect 298248 173023 298276 173051
rect 298310 173023 298338 173051
rect 298372 173023 298400 173051
rect 298434 173023 298462 173051
rect 298248 172961 298276 172989
rect 298310 172961 298338 172989
rect 298372 172961 298400 172989
rect 298434 172961 298462 172989
rect 298248 164147 298276 164175
rect 298310 164147 298338 164175
rect 298372 164147 298400 164175
rect 298434 164147 298462 164175
rect 298248 164085 298276 164113
rect 298310 164085 298338 164113
rect 298372 164085 298400 164113
rect 298434 164085 298462 164113
rect 298248 164023 298276 164051
rect 298310 164023 298338 164051
rect 298372 164023 298400 164051
rect 298434 164023 298462 164051
rect 298248 163961 298276 163989
rect 298310 163961 298338 163989
rect 298372 163961 298400 163989
rect 298434 163961 298462 163989
rect 298248 155147 298276 155175
rect 298310 155147 298338 155175
rect 298372 155147 298400 155175
rect 298434 155147 298462 155175
rect 298248 155085 298276 155113
rect 298310 155085 298338 155113
rect 298372 155085 298400 155113
rect 298434 155085 298462 155113
rect 298248 155023 298276 155051
rect 298310 155023 298338 155051
rect 298372 155023 298400 155051
rect 298434 155023 298462 155051
rect 298248 154961 298276 154989
rect 298310 154961 298338 154989
rect 298372 154961 298400 154989
rect 298434 154961 298462 154989
rect 298248 146147 298276 146175
rect 298310 146147 298338 146175
rect 298372 146147 298400 146175
rect 298434 146147 298462 146175
rect 298248 146085 298276 146113
rect 298310 146085 298338 146113
rect 298372 146085 298400 146113
rect 298434 146085 298462 146113
rect 298248 146023 298276 146051
rect 298310 146023 298338 146051
rect 298372 146023 298400 146051
rect 298434 146023 298462 146051
rect 298248 145961 298276 145989
rect 298310 145961 298338 145989
rect 298372 145961 298400 145989
rect 298434 145961 298462 145989
rect 298248 137147 298276 137175
rect 298310 137147 298338 137175
rect 298372 137147 298400 137175
rect 298434 137147 298462 137175
rect 298248 137085 298276 137113
rect 298310 137085 298338 137113
rect 298372 137085 298400 137113
rect 298434 137085 298462 137113
rect 298248 137023 298276 137051
rect 298310 137023 298338 137051
rect 298372 137023 298400 137051
rect 298434 137023 298462 137051
rect 298248 136961 298276 136989
rect 298310 136961 298338 136989
rect 298372 136961 298400 136989
rect 298434 136961 298462 136989
rect 298248 128147 298276 128175
rect 298310 128147 298338 128175
rect 298372 128147 298400 128175
rect 298434 128147 298462 128175
rect 298248 128085 298276 128113
rect 298310 128085 298338 128113
rect 298372 128085 298400 128113
rect 298434 128085 298462 128113
rect 298248 128023 298276 128051
rect 298310 128023 298338 128051
rect 298372 128023 298400 128051
rect 298434 128023 298462 128051
rect 298248 127961 298276 127989
rect 298310 127961 298338 127989
rect 298372 127961 298400 127989
rect 298434 127961 298462 127989
rect 298248 119147 298276 119175
rect 298310 119147 298338 119175
rect 298372 119147 298400 119175
rect 298434 119147 298462 119175
rect 298248 119085 298276 119113
rect 298310 119085 298338 119113
rect 298372 119085 298400 119113
rect 298434 119085 298462 119113
rect 298248 119023 298276 119051
rect 298310 119023 298338 119051
rect 298372 119023 298400 119051
rect 298434 119023 298462 119051
rect 298248 118961 298276 118989
rect 298310 118961 298338 118989
rect 298372 118961 298400 118989
rect 298434 118961 298462 118989
rect 298248 110147 298276 110175
rect 298310 110147 298338 110175
rect 298372 110147 298400 110175
rect 298434 110147 298462 110175
rect 298248 110085 298276 110113
rect 298310 110085 298338 110113
rect 298372 110085 298400 110113
rect 298434 110085 298462 110113
rect 298248 110023 298276 110051
rect 298310 110023 298338 110051
rect 298372 110023 298400 110051
rect 298434 110023 298462 110051
rect 298248 109961 298276 109989
rect 298310 109961 298338 109989
rect 298372 109961 298400 109989
rect 298434 109961 298462 109989
rect 298248 101147 298276 101175
rect 298310 101147 298338 101175
rect 298372 101147 298400 101175
rect 298434 101147 298462 101175
rect 298248 101085 298276 101113
rect 298310 101085 298338 101113
rect 298372 101085 298400 101113
rect 298434 101085 298462 101113
rect 298248 101023 298276 101051
rect 298310 101023 298338 101051
rect 298372 101023 298400 101051
rect 298434 101023 298462 101051
rect 298248 100961 298276 100989
rect 298310 100961 298338 100989
rect 298372 100961 298400 100989
rect 298434 100961 298462 100989
rect 298248 92147 298276 92175
rect 298310 92147 298338 92175
rect 298372 92147 298400 92175
rect 298434 92147 298462 92175
rect 298248 92085 298276 92113
rect 298310 92085 298338 92113
rect 298372 92085 298400 92113
rect 298434 92085 298462 92113
rect 298248 92023 298276 92051
rect 298310 92023 298338 92051
rect 298372 92023 298400 92051
rect 298434 92023 298462 92051
rect 298248 91961 298276 91989
rect 298310 91961 298338 91989
rect 298372 91961 298400 91989
rect 298434 91961 298462 91989
rect 298248 83147 298276 83175
rect 298310 83147 298338 83175
rect 298372 83147 298400 83175
rect 298434 83147 298462 83175
rect 298248 83085 298276 83113
rect 298310 83085 298338 83113
rect 298372 83085 298400 83113
rect 298434 83085 298462 83113
rect 298248 83023 298276 83051
rect 298310 83023 298338 83051
rect 298372 83023 298400 83051
rect 298434 83023 298462 83051
rect 298248 82961 298276 82989
rect 298310 82961 298338 82989
rect 298372 82961 298400 82989
rect 298434 82961 298462 82989
rect 298248 74147 298276 74175
rect 298310 74147 298338 74175
rect 298372 74147 298400 74175
rect 298434 74147 298462 74175
rect 298248 74085 298276 74113
rect 298310 74085 298338 74113
rect 298372 74085 298400 74113
rect 298434 74085 298462 74113
rect 298248 74023 298276 74051
rect 298310 74023 298338 74051
rect 298372 74023 298400 74051
rect 298434 74023 298462 74051
rect 298248 73961 298276 73989
rect 298310 73961 298338 73989
rect 298372 73961 298400 73989
rect 298434 73961 298462 73989
rect 298248 65147 298276 65175
rect 298310 65147 298338 65175
rect 298372 65147 298400 65175
rect 298434 65147 298462 65175
rect 298248 65085 298276 65113
rect 298310 65085 298338 65113
rect 298372 65085 298400 65113
rect 298434 65085 298462 65113
rect 298248 65023 298276 65051
rect 298310 65023 298338 65051
rect 298372 65023 298400 65051
rect 298434 65023 298462 65051
rect 298248 64961 298276 64989
rect 298310 64961 298338 64989
rect 298372 64961 298400 64989
rect 298434 64961 298462 64989
rect 298248 56147 298276 56175
rect 298310 56147 298338 56175
rect 298372 56147 298400 56175
rect 298434 56147 298462 56175
rect 298248 56085 298276 56113
rect 298310 56085 298338 56113
rect 298372 56085 298400 56113
rect 298434 56085 298462 56113
rect 298248 56023 298276 56051
rect 298310 56023 298338 56051
rect 298372 56023 298400 56051
rect 298434 56023 298462 56051
rect 298248 55961 298276 55989
rect 298310 55961 298338 55989
rect 298372 55961 298400 55989
rect 298434 55961 298462 55989
rect 298248 47147 298276 47175
rect 298310 47147 298338 47175
rect 298372 47147 298400 47175
rect 298434 47147 298462 47175
rect 298248 47085 298276 47113
rect 298310 47085 298338 47113
rect 298372 47085 298400 47113
rect 298434 47085 298462 47113
rect 298248 47023 298276 47051
rect 298310 47023 298338 47051
rect 298372 47023 298400 47051
rect 298434 47023 298462 47051
rect 298248 46961 298276 46989
rect 298310 46961 298338 46989
rect 298372 46961 298400 46989
rect 298434 46961 298462 46989
rect 298248 38147 298276 38175
rect 298310 38147 298338 38175
rect 298372 38147 298400 38175
rect 298434 38147 298462 38175
rect 298248 38085 298276 38113
rect 298310 38085 298338 38113
rect 298372 38085 298400 38113
rect 298434 38085 298462 38113
rect 298248 38023 298276 38051
rect 298310 38023 298338 38051
rect 298372 38023 298400 38051
rect 298434 38023 298462 38051
rect 298248 37961 298276 37989
rect 298310 37961 298338 37989
rect 298372 37961 298400 37989
rect 298434 37961 298462 37989
rect 298248 29147 298276 29175
rect 298310 29147 298338 29175
rect 298372 29147 298400 29175
rect 298434 29147 298462 29175
rect 298248 29085 298276 29113
rect 298310 29085 298338 29113
rect 298372 29085 298400 29113
rect 298434 29085 298462 29113
rect 298248 29023 298276 29051
rect 298310 29023 298338 29051
rect 298372 29023 298400 29051
rect 298434 29023 298462 29051
rect 298248 28961 298276 28989
rect 298310 28961 298338 28989
rect 298372 28961 298400 28989
rect 298434 28961 298462 28989
rect 298248 20147 298276 20175
rect 298310 20147 298338 20175
rect 298372 20147 298400 20175
rect 298434 20147 298462 20175
rect 298248 20085 298276 20113
rect 298310 20085 298338 20113
rect 298372 20085 298400 20113
rect 298434 20085 298462 20113
rect 298248 20023 298276 20051
rect 298310 20023 298338 20051
rect 298372 20023 298400 20051
rect 298434 20023 298462 20051
rect 298248 19961 298276 19989
rect 298310 19961 298338 19989
rect 298372 19961 298400 19989
rect 298434 19961 298462 19989
rect 298248 11147 298276 11175
rect 298310 11147 298338 11175
rect 298372 11147 298400 11175
rect 298434 11147 298462 11175
rect 298248 11085 298276 11113
rect 298310 11085 298338 11113
rect 298372 11085 298400 11113
rect 298434 11085 298462 11113
rect 298248 11023 298276 11051
rect 298310 11023 298338 11051
rect 298372 11023 298400 11051
rect 298434 11023 298462 11051
rect 298248 10961 298276 10989
rect 298310 10961 298338 10989
rect 298372 10961 298400 10989
rect 298434 10961 298462 10989
rect 298248 2147 298276 2175
rect 298310 2147 298338 2175
rect 298372 2147 298400 2175
rect 298434 2147 298462 2175
rect 298248 2085 298276 2113
rect 298310 2085 298338 2113
rect 298372 2085 298400 2113
rect 298434 2085 298462 2113
rect 298248 2023 298276 2051
rect 298310 2023 298338 2051
rect 298372 2023 298400 2051
rect 298434 2023 298462 2051
rect 298248 1961 298276 1989
rect 298310 1961 298338 1989
rect 298372 1961 298400 1989
rect 298434 1961 298462 1989
rect 298248 -108 298276 -80
rect 298310 -108 298338 -80
rect 298372 -108 298400 -80
rect 298434 -108 298462 -80
rect 298248 -170 298276 -142
rect 298310 -170 298338 -142
rect 298372 -170 298400 -142
rect 298434 -170 298462 -142
rect 298248 -232 298276 -204
rect 298310 -232 298338 -204
rect 298372 -232 298400 -204
rect 298434 -232 298462 -204
rect 298248 -294 298276 -266
rect 298310 -294 298338 -266
rect 298372 -294 298400 -266
rect 298434 -294 298462 -266
rect 298728 293147 298756 293175
rect 298790 293147 298818 293175
rect 298852 293147 298880 293175
rect 298914 293147 298942 293175
rect 298728 293085 298756 293113
rect 298790 293085 298818 293113
rect 298852 293085 298880 293113
rect 298914 293085 298942 293113
rect 298728 293023 298756 293051
rect 298790 293023 298818 293051
rect 298852 293023 298880 293051
rect 298914 293023 298942 293051
rect 298728 292961 298756 292989
rect 298790 292961 298818 292989
rect 298852 292961 298880 292989
rect 298914 292961 298942 292989
rect 298728 284147 298756 284175
rect 298790 284147 298818 284175
rect 298852 284147 298880 284175
rect 298914 284147 298942 284175
rect 298728 284085 298756 284113
rect 298790 284085 298818 284113
rect 298852 284085 298880 284113
rect 298914 284085 298942 284113
rect 298728 284023 298756 284051
rect 298790 284023 298818 284051
rect 298852 284023 298880 284051
rect 298914 284023 298942 284051
rect 298728 283961 298756 283989
rect 298790 283961 298818 283989
rect 298852 283961 298880 283989
rect 298914 283961 298942 283989
rect 298728 275147 298756 275175
rect 298790 275147 298818 275175
rect 298852 275147 298880 275175
rect 298914 275147 298942 275175
rect 298728 275085 298756 275113
rect 298790 275085 298818 275113
rect 298852 275085 298880 275113
rect 298914 275085 298942 275113
rect 298728 275023 298756 275051
rect 298790 275023 298818 275051
rect 298852 275023 298880 275051
rect 298914 275023 298942 275051
rect 298728 274961 298756 274989
rect 298790 274961 298818 274989
rect 298852 274961 298880 274989
rect 298914 274961 298942 274989
rect 298728 266147 298756 266175
rect 298790 266147 298818 266175
rect 298852 266147 298880 266175
rect 298914 266147 298942 266175
rect 298728 266085 298756 266113
rect 298790 266085 298818 266113
rect 298852 266085 298880 266113
rect 298914 266085 298942 266113
rect 298728 266023 298756 266051
rect 298790 266023 298818 266051
rect 298852 266023 298880 266051
rect 298914 266023 298942 266051
rect 298728 265961 298756 265989
rect 298790 265961 298818 265989
rect 298852 265961 298880 265989
rect 298914 265961 298942 265989
rect 298728 257147 298756 257175
rect 298790 257147 298818 257175
rect 298852 257147 298880 257175
rect 298914 257147 298942 257175
rect 298728 257085 298756 257113
rect 298790 257085 298818 257113
rect 298852 257085 298880 257113
rect 298914 257085 298942 257113
rect 298728 257023 298756 257051
rect 298790 257023 298818 257051
rect 298852 257023 298880 257051
rect 298914 257023 298942 257051
rect 298728 256961 298756 256989
rect 298790 256961 298818 256989
rect 298852 256961 298880 256989
rect 298914 256961 298942 256989
rect 298728 248147 298756 248175
rect 298790 248147 298818 248175
rect 298852 248147 298880 248175
rect 298914 248147 298942 248175
rect 298728 248085 298756 248113
rect 298790 248085 298818 248113
rect 298852 248085 298880 248113
rect 298914 248085 298942 248113
rect 298728 248023 298756 248051
rect 298790 248023 298818 248051
rect 298852 248023 298880 248051
rect 298914 248023 298942 248051
rect 298728 247961 298756 247989
rect 298790 247961 298818 247989
rect 298852 247961 298880 247989
rect 298914 247961 298942 247989
rect 298728 239147 298756 239175
rect 298790 239147 298818 239175
rect 298852 239147 298880 239175
rect 298914 239147 298942 239175
rect 298728 239085 298756 239113
rect 298790 239085 298818 239113
rect 298852 239085 298880 239113
rect 298914 239085 298942 239113
rect 298728 239023 298756 239051
rect 298790 239023 298818 239051
rect 298852 239023 298880 239051
rect 298914 239023 298942 239051
rect 298728 238961 298756 238989
rect 298790 238961 298818 238989
rect 298852 238961 298880 238989
rect 298914 238961 298942 238989
rect 298728 230147 298756 230175
rect 298790 230147 298818 230175
rect 298852 230147 298880 230175
rect 298914 230147 298942 230175
rect 298728 230085 298756 230113
rect 298790 230085 298818 230113
rect 298852 230085 298880 230113
rect 298914 230085 298942 230113
rect 298728 230023 298756 230051
rect 298790 230023 298818 230051
rect 298852 230023 298880 230051
rect 298914 230023 298942 230051
rect 298728 229961 298756 229989
rect 298790 229961 298818 229989
rect 298852 229961 298880 229989
rect 298914 229961 298942 229989
rect 298728 221147 298756 221175
rect 298790 221147 298818 221175
rect 298852 221147 298880 221175
rect 298914 221147 298942 221175
rect 298728 221085 298756 221113
rect 298790 221085 298818 221113
rect 298852 221085 298880 221113
rect 298914 221085 298942 221113
rect 298728 221023 298756 221051
rect 298790 221023 298818 221051
rect 298852 221023 298880 221051
rect 298914 221023 298942 221051
rect 298728 220961 298756 220989
rect 298790 220961 298818 220989
rect 298852 220961 298880 220989
rect 298914 220961 298942 220989
rect 298728 212147 298756 212175
rect 298790 212147 298818 212175
rect 298852 212147 298880 212175
rect 298914 212147 298942 212175
rect 298728 212085 298756 212113
rect 298790 212085 298818 212113
rect 298852 212085 298880 212113
rect 298914 212085 298942 212113
rect 298728 212023 298756 212051
rect 298790 212023 298818 212051
rect 298852 212023 298880 212051
rect 298914 212023 298942 212051
rect 298728 211961 298756 211989
rect 298790 211961 298818 211989
rect 298852 211961 298880 211989
rect 298914 211961 298942 211989
rect 298728 203147 298756 203175
rect 298790 203147 298818 203175
rect 298852 203147 298880 203175
rect 298914 203147 298942 203175
rect 298728 203085 298756 203113
rect 298790 203085 298818 203113
rect 298852 203085 298880 203113
rect 298914 203085 298942 203113
rect 298728 203023 298756 203051
rect 298790 203023 298818 203051
rect 298852 203023 298880 203051
rect 298914 203023 298942 203051
rect 298728 202961 298756 202989
rect 298790 202961 298818 202989
rect 298852 202961 298880 202989
rect 298914 202961 298942 202989
rect 298728 194147 298756 194175
rect 298790 194147 298818 194175
rect 298852 194147 298880 194175
rect 298914 194147 298942 194175
rect 298728 194085 298756 194113
rect 298790 194085 298818 194113
rect 298852 194085 298880 194113
rect 298914 194085 298942 194113
rect 298728 194023 298756 194051
rect 298790 194023 298818 194051
rect 298852 194023 298880 194051
rect 298914 194023 298942 194051
rect 298728 193961 298756 193989
rect 298790 193961 298818 193989
rect 298852 193961 298880 193989
rect 298914 193961 298942 193989
rect 298728 185147 298756 185175
rect 298790 185147 298818 185175
rect 298852 185147 298880 185175
rect 298914 185147 298942 185175
rect 298728 185085 298756 185113
rect 298790 185085 298818 185113
rect 298852 185085 298880 185113
rect 298914 185085 298942 185113
rect 298728 185023 298756 185051
rect 298790 185023 298818 185051
rect 298852 185023 298880 185051
rect 298914 185023 298942 185051
rect 298728 184961 298756 184989
rect 298790 184961 298818 184989
rect 298852 184961 298880 184989
rect 298914 184961 298942 184989
rect 298728 176147 298756 176175
rect 298790 176147 298818 176175
rect 298852 176147 298880 176175
rect 298914 176147 298942 176175
rect 298728 176085 298756 176113
rect 298790 176085 298818 176113
rect 298852 176085 298880 176113
rect 298914 176085 298942 176113
rect 298728 176023 298756 176051
rect 298790 176023 298818 176051
rect 298852 176023 298880 176051
rect 298914 176023 298942 176051
rect 298728 175961 298756 175989
rect 298790 175961 298818 175989
rect 298852 175961 298880 175989
rect 298914 175961 298942 175989
rect 298728 167147 298756 167175
rect 298790 167147 298818 167175
rect 298852 167147 298880 167175
rect 298914 167147 298942 167175
rect 298728 167085 298756 167113
rect 298790 167085 298818 167113
rect 298852 167085 298880 167113
rect 298914 167085 298942 167113
rect 298728 167023 298756 167051
rect 298790 167023 298818 167051
rect 298852 167023 298880 167051
rect 298914 167023 298942 167051
rect 298728 166961 298756 166989
rect 298790 166961 298818 166989
rect 298852 166961 298880 166989
rect 298914 166961 298942 166989
rect 298728 158147 298756 158175
rect 298790 158147 298818 158175
rect 298852 158147 298880 158175
rect 298914 158147 298942 158175
rect 298728 158085 298756 158113
rect 298790 158085 298818 158113
rect 298852 158085 298880 158113
rect 298914 158085 298942 158113
rect 298728 158023 298756 158051
rect 298790 158023 298818 158051
rect 298852 158023 298880 158051
rect 298914 158023 298942 158051
rect 298728 157961 298756 157989
rect 298790 157961 298818 157989
rect 298852 157961 298880 157989
rect 298914 157961 298942 157989
rect 298728 149147 298756 149175
rect 298790 149147 298818 149175
rect 298852 149147 298880 149175
rect 298914 149147 298942 149175
rect 298728 149085 298756 149113
rect 298790 149085 298818 149113
rect 298852 149085 298880 149113
rect 298914 149085 298942 149113
rect 298728 149023 298756 149051
rect 298790 149023 298818 149051
rect 298852 149023 298880 149051
rect 298914 149023 298942 149051
rect 298728 148961 298756 148989
rect 298790 148961 298818 148989
rect 298852 148961 298880 148989
rect 298914 148961 298942 148989
rect 298728 140147 298756 140175
rect 298790 140147 298818 140175
rect 298852 140147 298880 140175
rect 298914 140147 298942 140175
rect 298728 140085 298756 140113
rect 298790 140085 298818 140113
rect 298852 140085 298880 140113
rect 298914 140085 298942 140113
rect 298728 140023 298756 140051
rect 298790 140023 298818 140051
rect 298852 140023 298880 140051
rect 298914 140023 298942 140051
rect 298728 139961 298756 139989
rect 298790 139961 298818 139989
rect 298852 139961 298880 139989
rect 298914 139961 298942 139989
rect 298728 131147 298756 131175
rect 298790 131147 298818 131175
rect 298852 131147 298880 131175
rect 298914 131147 298942 131175
rect 298728 131085 298756 131113
rect 298790 131085 298818 131113
rect 298852 131085 298880 131113
rect 298914 131085 298942 131113
rect 298728 131023 298756 131051
rect 298790 131023 298818 131051
rect 298852 131023 298880 131051
rect 298914 131023 298942 131051
rect 298728 130961 298756 130989
rect 298790 130961 298818 130989
rect 298852 130961 298880 130989
rect 298914 130961 298942 130989
rect 298728 122147 298756 122175
rect 298790 122147 298818 122175
rect 298852 122147 298880 122175
rect 298914 122147 298942 122175
rect 298728 122085 298756 122113
rect 298790 122085 298818 122113
rect 298852 122085 298880 122113
rect 298914 122085 298942 122113
rect 298728 122023 298756 122051
rect 298790 122023 298818 122051
rect 298852 122023 298880 122051
rect 298914 122023 298942 122051
rect 298728 121961 298756 121989
rect 298790 121961 298818 121989
rect 298852 121961 298880 121989
rect 298914 121961 298942 121989
rect 298728 113147 298756 113175
rect 298790 113147 298818 113175
rect 298852 113147 298880 113175
rect 298914 113147 298942 113175
rect 298728 113085 298756 113113
rect 298790 113085 298818 113113
rect 298852 113085 298880 113113
rect 298914 113085 298942 113113
rect 298728 113023 298756 113051
rect 298790 113023 298818 113051
rect 298852 113023 298880 113051
rect 298914 113023 298942 113051
rect 298728 112961 298756 112989
rect 298790 112961 298818 112989
rect 298852 112961 298880 112989
rect 298914 112961 298942 112989
rect 298728 104147 298756 104175
rect 298790 104147 298818 104175
rect 298852 104147 298880 104175
rect 298914 104147 298942 104175
rect 298728 104085 298756 104113
rect 298790 104085 298818 104113
rect 298852 104085 298880 104113
rect 298914 104085 298942 104113
rect 298728 104023 298756 104051
rect 298790 104023 298818 104051
rect 298852 104023 298880 104051
rect 298914 104023 298942 104051
rect 298728 103961 298756 103989
rect 298790 103961 298818 103989
rect 298852 103961 298880 103989
rect 298914 103961 298942 103989
rect 298728 95147 298756 95175
rect 298790 95147 298818 95175
rect 298852 95147 298880 95175
rect 298914 95147 298942 95175
rect 298728 95085 298756 95113
rect 298790 95085 298818 95113
rect 298852 95085 298880 95113
rect 298914 95085 298942 95113
rect 298728 95023 298756 95051
rect 298790 95023 298818 95051
rect 298852 95023 298880 95051
rect 298914 95023 298942 95051
rect 298728 94961 298756 94989
rect 298790 94961 298818 94989
rect 298852 94961 298880 94989
rect 298914 94961 298942 94989
rect 298728 86147 298756 86175
rect 298790 86147 298818 86175
rect 298852 86147 298880 86175
rect 298914 86147 298942 86175
rect 298728 86085 298756 86113
rect 298790 86085 298818 86113
rect 298852 86085 298880 86113
rect 298914 86085 298942 86113
rect 298728 86023 298756 86051
rect 298790 86023 298818 86051
rect 298852 86023 298880 86051
rect 298914 86023 298942 86051
rect 298728 85961 298756 85989
rect 298790 85961 298818 85989
rect 298852 85961 298880 85989
rect 298914 85961 298942 85989
rect 298728 77147 298756 77175
rect 298790 77147 298818 77175
rect 298852 77147 298880 77175
rect 298914 77147 298942 77175
rect 298728 77085 298756 77113
rect 298790 77085 298818 77113
rect 298852 77085 298880 77113
rect 298914 77085 298942 77113
rect 298728 77023 298756 77051
rect 298790 77023 298818 77051
rect 298852 77023 298880 77051
rect 298914 77023 298942 77051
rect 298728 76961 298756 76989
rect 298790 76961 298818 76989
rect 298852 76961 298880 76989
rect 298914 76961 298942 76989
rect 298728 68147 298756 68175
rect 298790 68147 298818 68175
rect 298852 68147 298880 68175
rect 298914 68147 298942 68175
rect 298728 68085 298756 68113
rect 298790 68085 298818 68113
rect 298852 68085 298880 68113
rect 298914 68085 298942 68113
rect 298728 68023 298756 68051
rect 298790 68023 298818 68051
rect 298852 68023 298880 68051
rect 298914 68023 298942 68051
rect 298728 67961 298756 67989
rect 298790 67961 298818 67989
rect 298852 67961 298880 67989
rect 298914 67961 298942 67989
rect 298728 59147 298756 59175
rect 298790 59147 298818 59175
rect 298852 59147 298880 59175
rect 298914 59147 298942 59175
rect 298728 59085 298756 59113
rect 298790 59085 298818 59113
rect 298852 59085 298880 59113
rect 298914 59085 298942 59113
rect 298728 59023 298756 59051
rect 298790 59023 298818 59051
rect 298852 59023 298880 59051
rect 298914 59023 298942 59051
rect 298728 58961 298756 58989
rect 298790 58961 298818 58989
rect 298852 58961 298880 58989
rect 298914 58961 298942 58989
rect 298728 50147 298756 50175
rect 298790 50147 298818 50175
rect 298852 50147 298880 50175
rect 298914 50147 298942 50175
rect 298728 50085 298756 50113
rect 298790 50085 298818 50113
rect 298852 50085 298880 50113
rect 298914 50085 298942 50113
rect 298728 50023 298756 50051
rect 298790 50023 298818 50051
rect 298852 50023 298880 50051
rect 298914 50023 298942 50051
rect 298728 49961 298756 49989
rect 298790 49961 298818 49989
rect 298852 49961 298880 49989
rect 298914 49961 298942 49989
rect 298728 41147 298756 41175
rect 298790 41147 298818 41175
rect 298852 41147 298880 41175
rect 298914 41147 298942 41175
rect 298728 41085 298756 41113
rect 298790 41085 298818 41113
rect 298852 41085 298880 41113
rect 298914 41085 298942 41113
rect 298728 41023 298756 41051
rect 298790 41023 298818 41051
rect 298852 41023 298880 41051
rect 298914 41023 298942 41051
rect 298728 40961 298756 40989
rect 298790 40961 298818 40989
rect 298852 40961 298880 40989
rect 298914 40961 298942 40989
rect 298728 32147 298756 32175
rect 298790 32147 298818 32175
rect 298852 32147 298880 32175
rect 298914 32147 298942 32175
rect 298728 32085 298756 32113
rect 298790 32085 298818 32113
rect 298852 32085 298880 32113
rect 298914 32085 298942 32113
rect 298728 32023 298756 32051
rect 298790 32023 298818 32051
rect 298852 32023 298880 32051
rect 298914 32023 298942 32051
rect 298728 31961 298756 31989
rect 298790 31961 298818 31989
rect 298852 31961 298880 31989
rect 298914 31961 298942 31989
rect 298728 23147 298756 23175
rect 298790 23147 298818 23175
rect 298852 23147 298880 23175
rect 298914 23147 298942 23175
rect 298728 23085 298756 23113
rect 298790 23085 298818 23113
rect 298852 23085 298880 23113
rect 298914 23085 298942 23113
rect 298728 23023 298756 23051
rect 298790 23023 298818 23051
rect 298852 23023 298880 23051
rect 298914 23023 298942 23051
rect 298728 22961 298756 22989
rect 298790 22961 298818 22989
rect 298852 22961 298880 22989
rect 298914 22961 298942 22989
rect 298728 14147 298756 14175
rect 298790 14147 298818 14175
rect 298852 14147 298880 14175
rect 298914 14147 298942 14175
rect 298728 14085 298756 14113
rect 298790 14085 298818 14113
rect 298852 14085 298880 14113
rect 298914 14085 298942 14113
rect 298728 14023 298756 14051
rect 298790 14023 298818 14051
rect 298852 14023 298880 14051
rect 298914 14023 298942 14051
rect 298728 13961 298756 13989
rect 298790 13961 298818 13989
rect 298852 13961 298880 13989
rect 298914 13961 298942 13989
rect 298728 5147 298756 5175
rect 298790 5147 298818 5175
rect 298852 5147 298880 5175
rect 298914 5147 298942 5175
rect 298728 5085 298756 5113
rect 298790 5085 298818 5113
rect 298852 5085 298880 5113
rect 298914 5085 298942 5113
rect 298728 5023 298756 5051
rect 298790 5023 298818 5051
rect 298852 5023 298880 5051
rect 298914 5023 298942 5051
rect 298728 4961 298756 4989
rect 298790 4961 298818 4989
rect 298852 4961 298880 4989
rect 298914 4961 298942 4989
rect 296457 -588 296485 -560
rect 296519 -588 296547 -560
rect 296581 -588 296609 -560
rect 296643 -588 296671 -560
rect 296457 -650 296485 -622
rect 296519 -650 296547 -622
rect 296581 -650 296609 -622
rect 296643 -650 296671 -622
rect 296457 -712 296485 -684
rect 296519 -712 296547 -684
rect 296581 -712 296609 -684
rect 296643 -712 296671 -684
rect 296457 -774 296485 -746
rect 296519 -774 296547 -746
rect 296581 -774 296609 -746
rect 296643 -774 296671 -746
rect 298728 -588 298756 -560
rect 298790 -588 298818 -560
rect 298852 -588 298880 -560
rect 298914 -588 298942 -560
rect 298728 -650 298756 -622
rect 298790 -650 298818 -622
rect 298852 -650 298880 -622
rect 298914 -650 298942 -622
rect 298728 -712 298756 -684
rect 298790 -712 298818 -684
rect 298852 -712 298880 -684
rect 298914 -712 298942 -684
rect 298728 -774 298756 -746
rect 298790 -774 298818 -746
rect 298852 -774 298880 -746
rect 298914 -774 298942 -746
<< metal5 >>
rect -958 299086 298990 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect -958 299024 298990 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect -958 298962 298990 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect -958 298900 298990 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect -958 298824 298990 298872
rect -478 298606 298510 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect -478 298544 298510 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect -478 298482 298510 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect -478 298420 298510 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect -478 298344 298510 298392
rect -958 293175 298990 293223
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect -958 293113 298990 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect -958 293051 298990 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect -958 292989 298990 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect -958 292913 298990 292961
rect -958 290175 298990 290223
rect -958 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298990 290175
rect -958 290113 298990 290147
rect -958 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298990 290113
rect -958 290051 298990 290085
rect -958 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298990 290051
rect -958 289989 298990 290023
rect -958 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298990 289989
rect -958 289913 298990 289961
rect -958 284175 298990 284223
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect -958 284113 298990 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect -958 284051 298990 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect -958 283989 298990 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect -958 283913 298990 283961
rect -958 281175 298990 281223
rect -958 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298990 281175
rect -958 281113 298990 281147
rect -958 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298990 281113
rect -958 281051 298990 281085
rect -958 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298990 281051
rect -958 280989 298990 281023
rect -958 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298990 280989
rect -958 280913 298990 280961
rect -958 275175 298990 275223
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 109939 275175
rect 109967 275147 110001 275175
rect 110029 275147 125299 275175
rect 125327 275147 125361 275175
rect 125389 275147 140659 275175
rect 140687 275147 140721 275175
rect 140749 275147 156019 275175
rect 156047 275147 156081 275175
rect 156109 275147 171379 275175
rect 171407 275147 171441 275175
rect 171469 275147 186739 275175
rect 186767 275147 186801 275175
rect 186829 275147 202099 275175
rect 202127 275147 202161 275175
rect 202189 275147 217459 275175
rect 217487 275147 217521 275175
rect 217549 275147 232819 275175
rect 232847 275147 232881 275175
rect 232909 275147 248179 275175
rect 248207 275147 248241 275175
rect 248269 275147 263539 275175
rect 263567 275147 263601 275175
rect 263629 275147 278899 275175
rect 278927 275147 278961 275175
rect 278989 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect -958 275113 298990 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 109939 275113
rect 109967 275085 110001 275113
rect 110029 275085 125299 275113
rect 125327 275085 125361 275113
rect 125389 275085 140659 275113
rect 140687 275085 140721 275113
rect 140749 275085 156019 275113
rect 156047 275085 156081 275113
rect 156109 275085 171379 275113
rect 171407 275085 171441 275113
rect 171469 275085 186739 275113
rect 186767 275085 186801 275113
rect 186829 275085 202099 275113
rect 202127 275085 202161 275113
rect 202189 275085 217459 275113
rect 217487 275085 217521 275113
rect 217549 275085 232819 275113
rect 232847 275085 232881 275113
rect 232909 275085 248179 275113
rect 248207 275085 248241 275113
rect 248269 275085 263539 275113
rect 263567 275085 263601 275113
rect 263629 275085 278899 275113
rect 278927 275085 278961 275113
rect 278989 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect -958 275051 298990 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 109939 275051
rect 109967 275023 110001 275051
rect 110029 275023 125299 275051
rect 125327 275023 125361 275051
rect 125389 275023 140659 275051
rect 140687 275023 140721 275051
rect 140749 275023 156019 275051
rect 156047 275023 156081 275051
rect 156109 275023 171379 275051
rect 171407 275023 171441 275051
rect 171469 275023 186739 275051
rect 186767 275023 186801 275051
rect 186829 275023 202099 275051
rect 202127 275023 202161 275051
rect 202189 275023 217459 275051
rect 217487 275023 217521 275051
rect 217549 275023 232819 275051
rect 232847 275023 232881 275051
rect 232909 275023 248179 275051
rect 248207 275023 248241 275051
rect 248269 275023 263539 275051
rect 263567 275023 263601 275051
rect 263629 275023 278899 275051
rect 278927 275023 278961 275051
rect 278989 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect -958 274989 298990 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 109939 274989
rect 109967 274961 110001 274989
rect 110029 274961 125299 274989
rect 125327 274961 125361 274989
rect 125389 274961 140659 274989
rect 140687 274961 140721 274989
rect 140749 274961 156019 274989
rect 156047 274961 156081 274989
rect 156109 274961 171379 274989
rect 171407 274961 171441 274989
rect 171469 274961 186739 274989
rect 186767 274961 186801 274989
rect 186829 274961 202099 274989
rect 202127 274961 202161 274989
rect 202189 274961 217459 274989
rect 217487 274961 217521 274989
rect 217549 274961 232819 274989
rect 232847 274961 232881 274989
rect 232909 274961 248179 274989
rect 248207 274961 248241 274989
rect 248269 274961 263539 274989
rect 263567 274961 263601 274989
rect 263629 274961 278899 274989
rect 278927 274961 278961 274989
rect 278989 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect -958 274913 298990 274961
rect -958 272175 298990 272223
rect -958 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 102259 272175
rect 102287 272147 102321 272175
rect 102349 272147 117619 272175
rect 117647 272147 117681 272175
rect 117709 272147 132979 272175
rect 133007 272147 133041 272175
rect 133069 272147 148339 272175
rect 148367 272147 148401 272175
rect 148429 272147 163699 272175
rect 163727 272147 163761 272175
rect 163789 272147 179059 272175
rect 179087 272147 179121 272175
rect 179149 272147 194419 272175
rect 194447 272147 194481 272175
rect 194509 272147 209779 272175
rect 209807 272147 209841 272175
rect 209869 272147 225139 272175
rect 225167 272147 225201 272175
rect 225229 272147 240499 272175
rect 240527 272147 240561 272175
rect 240589 272147 255859 272175
rect 255887 272147 255921 272175
rect 255949 272147 271219 272175
rect 271247 272147 271281 272175
rect 271309 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298990 272175
rect -958 272113 298990 272147
rect -958 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 102259 272113
rect 102287 272085 102321 272113
rect 102349 272085 117619 272113
rect 117647 272085 117681 272113
rect 117709 272085 132979 272113
rect 133007 272085 133041 272113
rect 133069 272085 148339 272113
rect 148367 272085 148401 272113
rect 148429 272085 163699 272113
rect 163727 272085 163761 272113
rect 163789 272085 179059 272113
rect 179087 272085 179121 272113
rect 179149 272085 194419 272113
rect 194447 272085 194481 272113
rect 194509 272085 209779 272113
rect 209807 272085 209841 272113
rect 209869 272085 225139 272113
rect 225167 272085 225201 272113
rect 225229 272085 240499 272113
rect 240527 272085 240561 272113
rect 240589 272085 255859 272113
rect 255887 272085 255921 272113
rect 255949 272085 271219 272113
rect 271247 272085 271281 272113
rect 271309 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298990 272113
rect -958 272051 298990 272085
rect -958 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 102259 272051
rect 102287 272023 102321 272051
rect 102349 272023 117619 272051
rect 117647 272023 117681 272051
rect 117709 272023 132979 272051
rect 133007 272023 133041 272051
rect 133069 272023 148339 272051
rect 148367 272023 148401 272051
rect 148429 272023 163699 272051
rect 163727 272023 163761 272051
rect 163789 272023 179059 272051
rect 179087 272023 179121 272051
rect 179149 272023 194419 272051
rect 194447 272023 194481 272051
rect 194509 272023 209779 272051
rect 209807 272023 209841 272051
rect 209869 272023 225139 272051
rect 225167 272023 225201 272051
rect 225229 272023 240499 272051
rect 240527 272023 240561 272051
rect 240589 272023 255859 272051
rect 255887 272023 255921 272051
rect 255949 272023 271219 272051
rect 271247 272023 271281 272051
rect 271309 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298990 272051
rect -958 271989 298990 272023
rect -958 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 102259 271989
rect 102287 271961 102321 271989
rect 102349 271961 117619 271989
rect 117647 271961 117681 271989
rect 117709 271961 132979 271989
rect 133007 271961 133041 271989
rect 133069 271961 148339 271989
rect 148367 271961 148401 271989
rect 148429 271961 163699 271989
rect 163727 271961 163761 271989
rect 163789 271961 179059 271989
rect 179087 271961 179121 271989
rect 179149 271961 194419 271989
rect 194447 271961 194481 271989
rect 194509 271961 209779 271989
rect 209807 271961 209841 271989
rect 209869 271961 225139 271989
rect 225167 271961 225201 271989
rect 225229 271961 240499 271989
rect 240527 271961 240561 271989
rect 240589 271961 255859 271989
rect 255887 271961 255921 271989
rect 255949 271961 271219 271989
rect 271247 271961 271281 271989
rect 271309 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298990 271989
rect -958 271913 298990 271961
rect -958 266175 298990 266223
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 19977 266175
rect 20005 266147 20039 266175
rect 20067 266147 20101 266175
rect 20129 266147 20163 266175
rect 20191 266147 35337 266175
rect 35365 266147 35399 266175
rect 35427 266147 35461 266175
rect 35489 266147 35523 266175
rect 35551 266147 50697 266175
rect 50725 266147 50759 266175
rect 50787 266147 50821 266175
rect 50849 266147 50883 266175
rect 50911 266147 66057 266175
rect 66085 266147 66119 266175
rect 66147 266147 66181 266175
rect 66209 266147 66243 266175
rect 66271 266147 81417 266175
rect 81445 266147 81479 266175
rect 81507 266147 81541 266175
rect 81569 266147 81603 266175
rect 81631 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 109939 266175
rect 109967 266147 110001 266175
rect 110029 266147 125299 266175
rect 125327 266147 125361 266175
rect 125389 266147 140659 266175
rect 140687 266147 140721 266175
rect 140749 266147 156019 266175
rect 156047 266147 156081 266175
rect 156109 266147 171379 266175
rect 171407 266147 171441 266175
rect 171469 266147 186739 266175
rect 186767 266147 186801 266175
rect 186829 266147 202099 266175
rect 202127 266147 202161 266175
rect 202189 266147 217459 266175
rect 217487 266147 217521 266175
rect 217549 266147 232819 266175
rect 232847 266147 232881 266175
rect 232909 266147 248179 266175
rect 248207 266147 248241 266175
rect 248269 266147 263539 266175
rect 263567 266147 263601 266175
rect 263629 266147 278899 266175
rect 278927 266147 278961 266175
rect 278989 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect -958 266113 298990 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 19977 266113
rect 20005 266085 20039 266113
rect 20067 266085 20101 266113
rect 20129 266085 20163 266113
rect 20191 266085 35337 266113
rect 35365 266085 35399 266113
rect 35427 266085 35461 266113
rect 35489 266085 35523 266113
rect 35551 266085 50697 266113
rect 50725 266085 50759 266113
rect 50787 266085 50821 266113
rect 50849 266085 50883 266113
rect 50911 266085 66057 266113
rect 66085 266085 66119 266113
rect 66147 266085 66181 266113
rect 66209 266085 66243 266113
rect 66271 266085 81417 266113
rect 81445 266085 81479 266113
rect 81507 266085 81541 266113
rect 81569 266085 81603 266113
rect 81631 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 109939 266113
rect 109967 266085 110001 266113
rect 110029 266085 125299 266113
rect 125327 266085 125361 266113
rect 125389 266085 140659 266113
rect 140687 266085 140721 266113
rect 140749 266085 156019 266113
rect 156047 266085 156081 266113
rect 156109 266085 171379 266113
rect 171407 266085 171441 266113
rect 171469 266085 186739 266113
rect 186767 266085 186801 266113
rect 186829 266085 202099 266113
rect 202127 266085 202161 266113
rect 202189 266085 217459 266113
rect 217487 266085 217521 266113
rect 217549 266085 232819 266113
rect 232847 266085 232881 266113
rect 232909 266085 248179 266113
rect 248207 266085 248241 266113
rect 248269 266085 263539 266113
rect 263567 266085 263601 266113
rect 263629 266085 278899 266113
rect 278927 266085 278961 266113
rect 278989 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect -958 266051 298990 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 19977 266051
rect 20005 266023 20039 266051
rect 20067 266023 20101 266051
rect 20129 266023 20163 266051
rect 20191 266023 35337 266051
rect 35365 266023 35399 266051
rect 35427 266023 35461 266051
rect 35489 266023 35523 266051
rect 35551 266023 50697 266051
rect 50725 266023 50759 266051
rect 50787 266023 50821 266051
rect 50849 266023 50883 266051
rect 50911 266023 66057 266051
rect 66085 266023 66119 266051
rect 66147 266023 66181 266051
rect 66209 266023 66243 266051
rect 66271 266023 81417 266051
rect 81445 266023 81479 266051
rect 81507 266023 81541 266051
rect 81569 266023 81603 266051
rect 81631 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 109939 266051
rect 109967 266023 110001 266051
rect 110029 266023 125299 266051
rect 125327 266023 125361 266051
rect 125389 266023 140659 266051
rect 140687 266023 140721 266051
rect 140749 266023 156019 266051
rect 156047 266023 156081 266051
rect 156109 266023 171379 266051
rect 171407 266023 171441 266051
rect 171469 266023 186739 266051
rect 186767 266023 186801 266051
rect 186829 266023 202099 266051
rect 202127 266023 202161 266051
rect 202189 266023 217459 266051
rect 217487 266023 217521 266051
rect 217549 266023 232819 266051
rect 232847 266023 232881 266051
rect 232909 266023 248179 266051
rect 248207 266023 248241 266051
rect 248269 266023 263539 266051
rect 263567 266023 263601 266051
rect 263629 266023 278899 266051
rect 278927 266023 278961 266051
rect 278989 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect -958 265989 298990 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 19977 265989
rect 20005 265961 20039 265989
rect 20067 265961 20101 265989
rect 20129 265961 20163 265989
rect 20191 265961 35337 265989
rect 35365 265961 35399 265989
rect 35427 265961 35461 265989
rect 35489 265961 35523 265989
rect 35551 265961 50697 265989
rect 50725 265961 50759 265989
rect 50787 265961 50821 265989
rect 50849 265961 50883 265989
rect 50911 265961 66057 265989
rect 66085 265961 66119 265989
rect 66147 265961 66181 265989
rect 66209 265961 66243 265989
rect 66271 265961 81417 265989
rect 81445 265961 81479 265989
rect 81507 265961 81541 265989
rect 81569 265961 81603 265989
rect 81631 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 109939 265989
rect 109967 265961 110001 265989
rect 110029 265961 125299 265989
rect 125327 265961 125361 265989
rect 125389 265961 140659 265989
rect 140687 265961 140721 265989
rect 140749 265961 156019 265989
rect 156047 265961 156081 265989
rect 156109 265961 171379 265989
rect 171407 265961 171441 265989
rect 171469 265961 186739 265989
rect 186767 265961 186801 265989
rect 186829 265961 202099 265989
rect 202127 265961 202161 265989
rect 202189 265961 217459 265989
rect 217487 265961 217521 265989
rect 217549 265961 232819 265989
rect 232847 265961 232881 265989
rect 232909 265961 248179 265989
rect 248207 265961 248241 265989
rect 248269 265961 263539 265989
rect 263567 265961 263601 265989
rect 263629 265961 278899 265989
rect 278927 265961 278961 265989
rect 278989 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect -958 265913 298990 265961
rect -958 263175 298990 263223
rect -958 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 33477 263175
rect 33505 263147 33539 263175
rect 33567 263147 33601 263175
rect 33629 263147 33663 263175
rect 33691 263147 48837 263175
rect 48865 263147 48899 263175
rect 48927 263147 48961 263175
rect 48989 263147 49023 263175
rect 49051 263147 64197 263175
rect 64225 263147 64259 263175
rect 64287 263147 64321 263175
rect 64349 263147 64383 263175
rect 64411 263147 79557 263175
rect 79585 263147 79619 263175
rect 79647 263147 79681 263175
rect 79709 263147 79743 263175
rect 79771 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 102259 263175
rect 102287 263147 102321 263175
rect 102349 263147 117619 263175
rect 117647 263147 117681 263175
rect 117709 263147 132979 263175
rect 133007 263147 133041 263175
rect 133069 263147 148339 263175
rect 148367 263147 148401 263175
rect 148429 263147 163699 263175
rect 163727 263147 163761 263175
rect 163789 263147 179059 263175
rect 179087 263147 179121 263175
rect 179149 263147 194419 263175
rect 194447 263147 194481 263175
rect 194509 263147 209779 263175
rect 209807 263147 209841 263175
rect 209869 263147 225139 263175
rect 225167 263147 225201 263175
rect 225229 263147 240499 263175
rect 240527 263147 240561 263175
rect 240589 263147 255859 263175
rect 255887 263147 255921 263175
rect 255949 263147 271219 263175
rect 271247 263147 271281 263175
rect 271309 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298990 263175
rect -958 263113 298990 263147
rect -958 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 33477 263113
rect 33505 263085 33539 263113
rect 33567 263085 33601 263113
rect 33629 263085 33663 263113
rect 33691 263085 48837 263113
rect 48865 263085 48899 263113
rect 48927 263085 48961 263113
rect 48989 263085 49023 263113
rect 49051 263085 64197 263113
rect 64225 263085 64259 263113
rect 64287 263085 64321 263113
rect 64349 263085 64383 263113
rect 64411 263085 79557 263113
rect 79585 263085 79619 263113
rect 79647 263085 79681 263113
rect 79709 263085 79743 263113
rect 79771 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 102259 263113
rect 102287 263085 102321 263113
rect 102349 263085 117619 263113
rect 117647 263085 117681 263113
rect 117709 263085 132979 263113
rect 133007 263085 133041 263113
rect 133069 263085 148339 263113
rect 148367 263085 148401 263113
rect 148429 263085 163699 263113
rect 163727 263085 163761 263113
rect 163789 263085 179059 263113
rect 179087 263085 179121 263113
rect 179149 263085 194419 263113
rect 194447 263085 194481 263113
rect 194509 263085 209779 263113
rect 209807 263085 209841 263113
rect 209869 263085 225139 263113
rect 225167 263085 225201 263113
rect 225229 263085 240499 263113
rect 240527 263085 240561 263113
rect 240589 263085 255859 263113
rect 255887 263085 255921 263113
rect 255949 263085 271219 263113
rect 271247 263085 271281 263113
rect 271309 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298990 263113
rect -958 263051 298990 263085
rect -958 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 33477 263051
rect 33505 263023 33539 263051
rect 33567 263023 33601 263051
rect 33629 263023 33663 263051
rect 33691 263023 48837 263051
rect 48865 263023 48899 263051
rect 48927 263023 48961 263051
rect 48989 263023 49023 263051
rect 49051 263023 64197 263051
rect 64225 263023 64259 263051
rect 64287 263023 64321 263051
rect 64349 263023 64383 263051
rect 64411 263023 79557 263051
rect 79585 263023 79619 263051
rect 79647 263023 79681 263051
rect 79709 263023 79743 263051
rect 79771 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 102259 263051
rect 102287 263023 102321 263051
rect 102349 263023 117619 263051
rect 117647 263023 117681 263051
rect 117709 263023 132979 263051
rect 133007 263023 133041 263051
rect 133069 263023 148339 263051
rect 148367 263023 148401 263051
rect 148429 263023 163699 263051
rect 163727 263023 163761 263051
rect 163789 263023 179059 263051
rect 179087 263023 179121 263051
rect 179149 263023 194419 263051
rect 194447 263023 194481 263051
rect 194509 263023 209779 263051
rect 209807 263023 209841 263051
rect 209869 263023 225139 263051
rect 225167 263023 225201 263051
rect 225229 263023 240499 263051
rect 240527 263023 240561 263051
rect 240589 263023 255859 263051
rect 255887 263023 255921 263051
rect 255949 263023 271219 263051
rect 271247 263023 271281 263051
rect 271309 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298990 263051
rect -958 262989 298990 263023
rect -958 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 33477 262989
rect 33505 262961 33539 262989
rect 33567 262961 33601 262989
rect 33629 262961 33663 262989
rect 33691 262961 48837 262989
rect 48865 262961 48899 262989
rect 48927 262961 48961 262989
rect 48989 262961 49023 262989
rect 49051 262961 64197 262989
rect 64225 262961 64259 262989
rect 64287 262961 64321 262989
rect 64349 262961 64383 262989
rect 64411 262961 79557 262989
rect 79585 262961 79619 262989
rect 79647 262961 79681 262989
rect 79709 262961 79743 262989
rect 79771 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 102259 262989
rect 102287 262961 102321 262989
rect 102349 262961 117619 262989
rect 117647 262961 117681 262989
rect 117709 262961 132979 262989
rect 133007 262961 133041 262989
rect 133069 262961 148339 262989
rect 148367 262961 148401 262989
rect 148429 262961 163699 262989
rect 163727 262961 163761 262989
rect 163789 262961 179059 262989
rect 179087 262961 179121 262989
rect 179149 262961 194419 262989
rect 194447 262961 194481 262989
rect 194509 262961 209779 262989
rect 209807 262961 209841 262989
rect 209869 262961 225139 262989
rect 225167 262961 225201 262989
rect 225229 262961 240499 262989
rect 240527 262961 240561 262989
rect 240589 262961 255859 262989
rect 255887 262961 255921 262989
rect 255949 262961 271219 262989
rect 271247 262961 271281 262989
rect 271309 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298990 262989
rect -958 262913 298990 262961
rect -958 257175 298990 257223
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 19977 257175
rect 20005 257147 20039 257175
rect 20067 257147 20101 257175
rect 20129 257147 20163 257175
rect 20191 257147 35337 257175
rect 35365 257147 35399 257175
rect 35427 257147 35461 257175
rect 35489 257147 35523 257175
rect 35551 257147 50697 257175
rect 50725 257147 50759 257175
rect 50787 257147 50821 257175
rect 50849 257147 50883 257175
rect 50911 257147 66057 257175
rect 66085 257147 66119 257175
rect 66147 257147 66181 257175
rect 66209 257147 66243 257175
rect 66271 257147 81417 257175
rect 81445 257147 81479 257175
rect 81507 257147 81541 257175
rect 81569 257147 81603 257175
rect 81631 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 109939 257175
rect 109967 257147 110001 257175
rect 110029 257147 125299 257175
rect 125327 257147 125361 257175
rect 125389 257147 140659 257175
rect 140687 257147 140721 257175
rect 140749 257147 156019 257175
rect 156047 257147 156081 257175
rect 156109 257147 171379 257175
rect 171407 257147 171441 257175
rect 171469 257147 186739 257175
rect 186767 257147 186801 257175
rect 186829 257147 202099 257175
rect 202127 257147 202161 257175
rect 202189 257147 217459 257175
rect 217487 257147 217521 257175
rect 217549 257147 232819 257175
rect 232847 257147 232881 257175
rect 232909 257147 248179 257175
rect 248207 257147 248241 257175
rect 248269 257147 263539 257175
rect 263567 257147 263601 257175
rect 263629 257147 278899 257175
rect 278927 257147 278961 257175
rect 278989 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect -958 257113 298990 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 19977 257113
rect 20005 257085 20039 257113
rect 20067 257085 20101 257113
rect 20129 257085 20163 257113
rect 20191 257085 35337 257113
rect 35365 257085 35399 257113
rect 35427 257085 35461 257113
rect 35489 257085 35523 257113
rect 35551 257085 50697 257113
rect 50725 257085 50759 257113
rect 50787 257085 50821 257113
rect 50849 257085 50883 257113
rect 50911 257085 66057 257113
rect 66085 257085 66119 257113
rect 66147 257085 66181 257113
rect 66209 257085 66243 257113
rect 66271 257085 81417 257113
rect 81445 257085 81479 257113
rect 81507 257085 81541 257113
rect 81569 257085 81603 257113
rect 81631 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 109939 257113
rect 109967 257085 110001 257113
rect 110029 257085 125299 257113
rect 125327 257085 125361 257113
rect 125389 257085 140659 257113
rect 140687 257085 140721 257113
rect 140749 257085 156019 257113
rect 156047 257085 156081 257113
rect 156109 257085 171379 257113
rect 171407 257085 171441 257113
rect 171469 257085 186739 257113
rect 186767 257085 186801 257113
rect 186829 257085 202099 257113
rect 202127 257085 202161 257113
rect 202189 257085 217459 257113
rect 217487 257085 217521 257113
rect 217549 257085 232819 257113
rect 232847 257085 232881 257113
rect 232909 257085 248179 257113
rect 248207 257085 248241 257113
rect 248269 257085 263539 257113
rect 263567 257085 263601 257113
rect 263629 257085 278899 257113
rect 278927 257085 278961 257113
rect 278989 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect -958 257051 298990 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 19977 257051
rect 20005 257023 20039 257051
rect 20067 257023 20101 257051
rect 20129 257023 20163 257051
rect 20191 257023 35337 257051
rect 35365 257023 35399 257051
rect 35427 257023 35461 257051
rect 35489 257023 35523 257051
rect 35551 257023 50697 257051
rect 50725 257023 50759 257051
rect 50787 257023 50821 257051
rect 50849 257023 50883 257051
rect 50911 257023 66057 257051
rect 66085 257023 66119 257051
rect 66147 257023 66181 257051
rect 66209 257023 66243 257051
rect 66271 257023 81417 257051
rect 81445 257023 81479 257051
rect 81507 257023 81541 257051
rect 81569 257023 81603 257051
rect 81631 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 109939 257051
rect 109967 257023 110001 257051
rect 110029 257023 125299 257051
rect 125327 257023 125361 257051
rect 125389 257023 140659 257051
rect 140687 257023 140721 257051
rect 140749 257023 156019 257051
rect 156047 257023 156081 257051
rect 156109 257023 171379 257051
rect 171407 257023 171441 257051
rect 171469 257023 186739 257051
rect 186767 257023 186801 257051
rect 186829 257023 202099 257051
rect 202127 257023 202161 257051
rect 202189 257023 217459 257051
rect 217487 257023 217521 257051
rect 217549 257023 232819 257051
rect 232847 257023 232881 257051
rect 232909 257023 248179 257051
rect 248207 257023 248241 257051
rect 248269 257023 263539 257051
rect 263567 257023 263601 257051
rect 263629 257023 278899 257051
rect 278927 257023 278961 257051
rect 278989 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect -958 256989 298990 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 19977 256989
rect 20005 256961 20039 256989
rect 20067 256961 20101 256989
rect 20129 256961 20163 256989
rect 20191 256961 35337 256989
rect 35365 256961 35399 256989
rect 35427 256961 35461 256989
rect 35489 256961 35523 256989
rect 35551 256961 50697 256989
rect 50725 256961 50759 256989
rect 50787 256961 50821 256989
rect 50849 256961 50883 256989
rect 50911 256961 66057 256989
rect 66085 256961 66119 256989
rect 66147 256961 66181 256989
rect 66209 256961 66243 256989
rect 66271 256961 81417 256989
rect 81445 256961 81479 256989
rect 81507 256961 81541 256989
rect 81569 256961 81603 256989
rect 81631 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 109939 256989
rect 109967 256961 110001 256989
rect 110029 256961 125299 256989
rect 125327 256961 125361 256989
rect 125389 256961 140659 256989
rect 140687 256961 140721 256989
rect 140749 256961 156019 256989
rect 156047 256961 156081 256989
rect 156109 256961 171379 256989
rect 171407 256961 171441 256989
rect 171469 256961 186739 256989
rect 186767 256961 186801 256989
rect 186829 256961 202099 256989
rect 202127 256961 202161 256989
rect 202189 256961 217459 256989
rect 217487 256961 217521 256989
rect 217549 256961 232819 256989
rect 232847 256961 232881 256989
rect 232909 256961 248179 256989
rect 248207 256961 248241 256989
rect 248269 256961 263539 256989
rect 263567 256961 263601 256989
rect 263629 256961 278899 256989
rect 278927 256961 278961 256989
rect 278989 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect -958 256913 298990 256961
rect -958 254175 298990 254223
rect -958 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 33477 254175
rect 33505 254147 33539 254175
rect 33567 254147 33601 254175
rect 33629 254147 33663 254175
rect 33691 254147 48837 254175
rect 48865 254147 48899 254175
rect 48927 254147 48961 254175
rect 48989 254147 49023 254175
rect 49051 254147 64197 254175
rect 64225 254147 64259 254175
rect 64287 254147 64321 254175
rect 64349 254147 64383 254175
rect 64411 254147 79557 254175
rect 79585 254147 79619 254175
rect 79647 254147 79681 254175
rect 79709 254147 79743 254175
rect 79771 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 102259 254175
rect 102287 254147 102321 254175
rect 102349 254147 117619 254175
rect 117647 254147 117681 254175
rect 117709 254147 132979 254175
rect 133007 254147 133041 254175
rect 133069 254147 148339 254175
rect 148367 254147 148401 254175
rect 148429 254147 163699 254175
rect 163727 254147 163761 254175
rect 163789 254147 179059 254175
rect 179087 254147 179121 254175
rect 179149 254147 194419 254175
rect 194447 254147 194481 254175
rect 194509 254147 209779 254175
rect 209807 254147 209841 254175
rect 209869 254147 225139 254175
rect 225167 254147 225201 254175
rect 225229 254147 240499 254175
rect 240527 254147 240561 254175
rect 240589 254147 255859 254175
rect 255887 254147 255921 254175
rect 255949 254147 271219 254175
rect 271247 254147 271281 254175
rect 271309 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298990 254175
rect -958 254113 298990 254147
rect -958 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 33477 254113
rect 33505 254085 33539 254113
rect 33567 254085 33601 254113
rect 33629 254085 33663 254113
rect 33691 254085 48837 254113
rect 48865 254085 48899 254113
rect 48927 254085 48961 254113
rect 48989 254085 49023 254113
rect 49051 254085 64197 254113
rect 64225 254085 64259 254113
rect 64287 254085 64321 254113
rect 64349 254085 64383 254113
rect 64411 254085 79557 254113
rect 79585 254085 79619 254113
rect 79647 254085 79681 254113
rect 79709 254085 79743 254113
rect 79771 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 102259 254113
rect 102287 254085 102321 254113
rect 102349 254085 117619 254113
rect 117647 254085 117681 254113
rect 117709 254085 132979 254113
rect 133007 254085 133041 254113
rect 133069 254085 148339 254113
rect 148367 254085 148401 254113
rect 148429 254085 163699 254113
rect 163727 254085 163761 254113
rect 163789 254085 179059 254113
rect 179087 254085 179121 254113
rect 179149 254085 194419 254113
rect 194447 254085 194481 254113
rect 194509 254085 209779 254113
rect 209807 254085 209841 254113
rect 209869 254085 225139 254113
rect 225167 254085 225201 254113
rect 225229 254085 240499 254113
rect 240527 254085 240561 254113
rect 240589 254085 255859 254113
rect 255887 254085 255921 254113
rect 255949 254085 271219 254113
rect 271247 254085 271281 254113
rect 271309 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298990 254113
rect -958 254051 298990 254085
rect -958 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 33477 254051
rect 33505 254023 33539 254051
rect 33567 254023 33601 254051
rect 33629 254023 33663 254051
rect 33691 254023 48837 254051
rect 48865 254023 48899 254051
rect 48927 254023 48961 254051
rect 48989 254023 49023 254051
rect 49051 254023 64197 254051
rect 64225 254023 64259 254051
rect 64287 254023 64321 254051
rect 64349 254023 64383 254051
rect 64411 254023 79557 254051
rect 79585 254023 79619 254051
rect 79647 254023 79681 254051
rect 79709 254023 79743 254051
rect 79771 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 102259 254051
rect 102287 254023 102321 254051
rect 102349 254023 117619 254051
rect 117647 254023 117681 254051
rect 117709 254023 132979 254051
rect 133007 254023 133041 254051
rect 133069 254023 148339 254051
rect 148367 254023 148401 254051
rect 148429 254023 163699 254051
rect 163727 254023 163761 254051
rect 163789 254023 179059 254051
rect 179087 254023 179121 254051
rect 179149 254023 194419 254051
rect 194447 254023 194481 254051
rect 194509 254023 209779 254051
rect 209807 254023 209841 254051
rect 209869 254023 225139 254051
rect 225167 254023 225201 254051
rect 225229 254023 240499 254051
rect 240527 254023 240561 254051
rect 240589 254023 255859 254051
rect 255887 254023 255921 254051
rect 255949 254023 271219 254051
rect 271247 254023 271281 254051
rect 271309 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298990 254051
rect -958 253989 298990 254023
rect -958 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 33477 253989
rect 33505 253961 33539 253989
rect 33567 253961 33601 253989
rect 33629 253961 33663 253989
rect 33691 253961 48837 253989
rect 48865 253961 48899 253989
rect 48927 253961 48961 253989
rect 48989 253961 49023 253989
rect 49051 253961 64197 253989
rect 64225 253961 64259 253989
rect 64287 253961 64321 253989
rect 64349 253961 64383 253989
rect 64411 253961 79557 253989
rect 79585 253961 79619 253989
rect 79647 253961 79681 253989
rect 79709 253961 79743 253989
rect 79771 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 102259 253989
rect 102287 253961 102321 253989
rect 102349 253961 117619 253989
rect 117647 253961 117681 253989
rect 117709 253961 132979 253989
rect 133007 253961 133041 253989
rect 133069 253961 148339 253989
rect 148367 253961 148401 253989
rect 148429 253961 163699 253989
rect 163727 253961 163761 253989
rect 163789 253961 179059 253989
rect 179087 253961 179121 253989
rect 179149 253961 194419 253989
rect 194447 253961 194481 253989
rect 194509 253961 209779 253989
rect 209807 253961 209841 253989
rect 209869 253961 225139 253989
rect 225167 253961 225201 253989
rect 225229 253961 240499 253989
rect 240527 253961 240561 253989
rect 240589 253961 255859 253989
rect 255887 253961 255921 253989
rect 255949 253961 271219 253989
rect 271247 253961 271281 253989
rect 271309 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298990 253989
rect -958 253913 298990 253961
rect -958 248175 298990 248223
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 19977 248175
rect 20005 248147 20039 248175
rect 20067 248147 20101 248175
rect 20129 248147 20163 248175
rect 20191 248147 35337 248175
rect 35365 248147 35399 248175
rect 35427 248147 35461 248175
rect 35489 248147 35523 248175
rect 35551 248147 50697 248175
rect 50725 248147 50759 248175
rect 50787 248147 50821 248175
rect 50849 248147 50883 248175
rect 50911 248147 66057 248175
rect 66085 248147 66119 248175
rect 66147 248147 66181 248175
rect 66209 248147 66243 248175
rect 66271 248147 81417 248175
rect 81445 248147 81479 248175
rect 81507 248147 81541 248175
rect 81569 248147 81603 248175
rect 81631 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 109939 248175
rect 109967 248147 110001 248175
rect 110029 248147 125299 248175
rect 125327 248147 125361 248175
rect 125389 248147 140659 248175
rect 140687 248147 140721 248175
rect 140749 248147 156019 248175
rect 156047 248147 156081 248175
rect 156109 248147 171379 248175
rect 171407 248147 171441 248175
rect 171469 248147 186739 248175
rect 186767 248147 186801 248175
rect 186829 248147 202099 248175
rect 202127 248147 202161 248175
rect 202189 248147 217459 248175
rect 217487 248147 217521 248175
rect 217549 248147 232819 248175
rect 232847 248147 232881 248175
rect 232909 248147 248179 248175
rect 248207 248147 248241 248175
rect 248269 248147 263539 248175
rect 263567 248147 263601 248175
rect 263629 248147 278899 248175
rect 278927 248147 278961 248175
rect 278989 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect -958 248113 298990 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 19977 248113
rect 20005 248085 20039 248113
rect 20067 248085 20101 248113
rect 20129 248085 20163 248113
rect 20191 248085 35337 248113
rect 35365 248085 35399 248113
rect 35427 248085 35461 248113
rect 35489 248085 35523 248113
rect 35551 248085 50697 248113
rect 50725 248085 50759 248113
rect 50787 248085 50821 248113
rect 50849 248085 50883 248113
rect 50911 248085 66057 248113
rect 66085 248085 66119 248113
rect 66147 248085 66181 248113
rect 66209 248085 66243 248113
rect 66271 248085 81417 248113
rect 81445 248085 81479 248113
rect 81507 248085 81541 248113
rect 81569 248085 81603 248113
rect 81631 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 109939 248113
rect 109967 248085 110001 248113
rect 110029 248085 125299 248113
rect 125327 248085 125361 248113
rect 125389 248085 140659 248113
rect 140687 248085 140721 248113
rect 140749 248085 156019 248113
rect 156047 248085 156081 248113
rect 156109 248085 171379 248113
rect 171407 248085 171441 248113
rect 171469 248085 186739 248113
rect 186767 248085 186801 248113
rect 186829 248085 202099 248113
rect 202127 248085 202161 248113
rect 202189 248085 217459 248113
rect 217487 248085 217521 248113
rect 217549 248085 232819 248113
rect 232847 248085 232881 248113
rect 232909 248085 248179 248113
rect 248207 248085 248241 248113
rect 248269 248085 263539 248113
rect 263567 248085 263601 248113
rect 263629 248085 278899 248113
rect 278927 248085 278961 248113
rect 278989 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect -958 248051 298990 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 19977 248051
rect 20005 248023 20039 248051
rect 20067 248023 20101 248051
rect 20129 248023 20163 248051
rect 20191 248023 35337 248051
rect 35365 248023 35399 248051
rect 35427 248023 35461 248051
rect 35489 248023 35523 248051
rect 35551 248023 50697 248051
rect 50725 248023 50759 248051
rect 50787 248023 50821 248051
rect 50849 248023 50883 248051
rect 50911 248023 66057 248051
rect 66085 248023 66119 248051
rect 66147 248023 66181 248051
rect 66209 248023 66243 248051
rect 66271 248023 81417 248051
rect 81445 248023 81479 248051
rect 81507 248023 81541 248051
rect 81569 248023 81603 248051
rect 81631 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 109939 248051
rect 109967 248023 110001 248051
rect 110029 248023 125299 248051
rect 125327 248023 125361 248051
rect 125389 248023 140659 248051
rect 140687 248023 140721 248051
rect 140749 248023 156019 248051
rect 156047 248023 156081 248051
rect 156109 248023 171379 248051
rect 171407 248023 171441 248051
rect 171469 248023 186739 248051
rect 186767 248023 186801 248051
rect 186829 248023 202099 248051
rect 202127 248023 202161 248051
rect 202189 248023 217459 248051
rect 217487 248023 217521 248051
rect 217549 248023 232819 248051
rect 232847 248023 232881 248051
rect 232909 248023 248179 248051
rect 248207 248023 248241 248051
rect 248269 248023 263539 248051
rect 263567 248023 263601 248051
rect 263629 248023 278899 248051
rect 278927 248023 278961 248051
rect 278989 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect -958 247989 298990 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 19977 247989
rect 20005 247961 20039 247989
rect 20067 247961 20101 247989
rect 20129 247961 20163 247989
rect 20191 247961 35337 247989
rect 35365 247961 35399 247989
rect 35427 247961 35461 247989
rect 35489 247961 35523 247989
rect 35551 247961 50697 247989
rect 50725 247961 50759 247989
rect 50787 247961 50821 247989
rect 50849 247961 50883 247989
rect 50911 247961 66057 247989
rect 66085 247961 66119 247989
rect 66147 247961 66181 247989
rect 66209 247961 66243 247989
rect 66271 247961 81417 247989
rect 81445 247961 81479 247989
rect 81507 247961 81541 247989
rect 81569 247961 81603 247989
rect 81631 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 109939 247989
rect 109967 247961 110001 247989
rect 110029 247961 125299 247989
rect 125327 247961 125361 247989
rect 125389 247961 140659 247989
rect 140687 247961 140721 247989
rect 140749 247961 156019 247989
rect 156047 247961 156081 247989
rect 156109 247961 171379 247989
rect 171407 247961 171441 247989
rect 171469 247961 186739 247989
rect 186767 247961 186801 247989
rect 186829 247961 202099 247989
rect 202127 247961 202161 247989
rect 202189 247961 217459 247989
rect 217487 247961 217521 247989
rect 217549 247961 232819 247989
rect 232847 247961 232881 247989
rect 232909 247961 248179 247989
rect 248207 247961 248241 247989
rect 248269 247961 263539 247989
rect 263567 247961 263601 247989
rect 263629 247961 278899 247989
rect 278927 247961 278961 247989
rect 278989 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect -958 247913 298990 247961
rect -958 245175 298990 245223
rect -958 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 33477 245175
rect 33505 245147 33539 245175
rect 33567 245147 33601 245175
rect 33629 245147 33663 245175
rect 33691 245147 48837 245175
rect 48865 245147 48899 245175
rect 48927 245147 48961 245175
rect 48989 245147 49023 245175
rect 49051 245147 64197 245175
rect 64225 245147 64259 245175
rect 64287 245147 64321 245175
rect 64349 245147 64383 245175
rect 64411 245147 79557 245175
rect 79585 245147 79619 245175
rect 79647 245147 79681 245175
rect 79709 245147 79743 245175
rect 79771 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 102259 245175
rect 102287 245147 102321 245175
rect 102349 245147 117619 245175
rect 117647 245147 117681 245175
rect 117709 245147 132979 245175
rect 133007 245147 133041 245175
rect 133069 245147 148339 245175
rect 148367 245147 148401 245175
rect 148429 245147 163699 245175
rect 163727 245147 163761 245175
rect 163789 245147 179059 245175
rect 179087 245147 179121 245175
rect 179149 245147 194419 245175
rect 194447 245147 194481 245175
rect 194509 245147 209779 245175
rect 209807 245147 209841 245175
rect 209869 245147 225139 245175
rect 225167 245147 225201 245175
rect 225229 245147 240499 245175
rect 240527 245147 240561 245175
rect 240589 245147 255859 245175
rect 255887 245147 255921 245175
rect 255949 245147 271219 245175
rect 271247 245147 271281 245175
rect 271309 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298990 245175
rect -958 245113 298990 245147
rect -958 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 33477 245113
rect 33505 245085 33539 245113
rect 33567 245085 33601 245113
rect 33629 245085 33663 245113
rect 33691 245085 48837 245113
rect 48865 245085 48899 245113
rect 48927 245085 48961 245113
rect 48989 245085 49023 245113
rect 49051 245085 64197 245113
rect 64225 245085 64259 245113
rect 64287 245085 64321 245113
rect 64349 245085 64383 245113
rect 64411 245085 79557 245113
rect 79585 245085 79619 245113
rect 79647 245085 79681 245113
rect 79709 245085 79743 245113
rect 79771 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 102259 245113
rect 102287 245085 102321 245113
rect 102349 245085 117619 245113
rect 117647 245085 117681 245113
rect 117709 245085 132979 245113
rect 133007 245085 133041 245113
rect 133069 245085 148339 245113
rect 148367 245085 148401 245113
rect 148429 245085 163699 245113
rect 163727 245085 163761 245113
rect 163789 245085 179059 245113
rect 179087 245085 179121 245113
rect 179149 245085 194419 245113
rect 194447 245085 194481 245113
rect 194509 245085 209779 245113
rect 209807 245085 209841 245113
rect 209869 245085 225139 245113
rect 225167 245085 225201 245113
rect 225229 245085 240499 245113
rect 240527 245085 240561 245113
rect 240589 245085 255859 245113
rect 255887 245085 255921 245113
rect 255949 245085 271219 245113
rect 271247 245085 271281 245113
rect 271309 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298990 245113
rect -958 245051 298990 245085
rect -958 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 33477 245051
rect 33505 245023 33539 245051
rect 33567 245023 33601 245051
rect 33629 245023 33663 245051
rect 33691 245023 48837 245051
rect 48865 245023 48899 245051
rect 48927 245023 48961 245051
rect 48989 245023 49023 245051
rect 49051 245023 64197 245051
rect 64225 245023 64259 245051
rect 64287 245023 64321 245051
rect 64349 245023 64383 245051
rect 64411 245023 79557 245051
rect 79585 245023 79619 245051
rect 79647 245023 79681 245051
rect 79709 245023 79743 245051
rect 79771 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 102259 245051
rect 102287 245023 102321 245051
rect 102349 245023 117619 245051
rect 117647 245023 117681 245051
rect 117709 245023 132979 245051
rect 133007 245023 133041 245051
rect 133069 245023 148339 245051
rect 148367 245023 148401 245051
rect 148429 245023 163699 245051
rect 163727 245023 163761 245051
rect 163789 245023 179059 245051
rect 179087 245023 179121 245051
rect 179149 245023 194419 245051
rect 194447 245023 194481 245051
rect 194509 245023 209779 245051
rect 209807 245023 209841 245051
rect 209869 245023 225139 245051
rect 225167 245023 225201 245051
rect 225229 245023 240499 245051
rect 240527 245023 240561 245051
rect 240589 245023 255859 245051
rect 255887 245023 255921 245051
rect 255949 245023 271219 245051
rect 271247 245023 271281 245051
rect 271309 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298990 245051
rect -958 244989 298990 245023
rect -958 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 33477 244989
rect 33505 244961 33539 244989
rect 33567 244961 33601 244989
rect 33629 244961 33663 244989
rect 33691 244961 48837 244989
rect 48865 244961 48899 244989
rect 48927 244961 48961 244989
rect 48989 244961 49023 244989
rect 49051 244961 64197 244989
rect 64225 244961 64259 244989
rect 64287 244961 64321 244989
rect 64349 244961 64383 244989
rect 64411 244961 79557 244989
rect 79585 244961 79619 244989
rect 79647 244961 79681 244989
rect 79709 244961 79743 244989
rect 79771 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 102259 244989
rect 102287 244961 102321 244989
rect 102349 244961 117619 244989
rect 117647 244961 117681 244989
rect 117709 244961 132979 244989
rect 133007 244961 133041 244989
rect 133069 244961 148339 244989
rect 148367 244961 148401 244989
rect 148429 244961 163699 244989
rect 163727 244961 163761 244989
rect 163789 244961 179059 244989
rect 179087 244961 179121 244989
rect 179149 244961 194419 244989
rect 194447 244961 194481 244989
rect 194509 244961 209779 244989
rect 209807 244961 209841 244989
rect 209869 244961 225139 244989
rect 225167 244961 225201 244989
rect 225229 244961 240499 244989
rect 240527 244961 240561 244989
rect 240589 244961 255859 244989
rect 255887 244961 255921 244989
rect 255949 244961 271219 244989
rect 271247 244961 271281 244989
rect 271309 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298990 244989
rect -958 244913 298990 244961
rect -958 239175 298990 239223
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 19977 239175
rect 20005 239147 20039 239175
rect 20067 239147 20101 239175
rect 20129 239147 20163 239175
rect 20191 239147 35337 239175
rect 35365 239147 35399 239175
rect 35427 239147 35461 239175
rect 35489 239147 35523 239175
rect 35551 239147 50697 239175
rect 50725 239147 50759 239175
rect 50787 239147 50821 239175
rect 50849 239147 50883 239175
rect 50911 239147 66057 239175
rect 66085 239147 66119 239175
rect 66147 239147 66181 239175
rect 66209 239147 66243 239175
rect 66271 239147 81417 239175
rect 81445 239147 81479 239175
rect 81507 239147 81541 239175
rect 81569 239147 81603 239175
rect 81631 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 109939 239175
rect 109967 239147 110001 239175
rect 110029 239147 125299 239175
rect 125327 239147 125361 239175
rect 125389 239147 140659 239175
rect 140687 239147 140721 239175
rect 140749 239147 156019 239175
rect 156047 239147 156081 239175
rect 156109 239147 171379 239175
rect 171407 239147 171441 239175
rect 171469 239147 186739 239175
rect 186767 239147 186801 239175
rect 186829 239147 202099 239175
rect 202127 239147 202161 239175
rect 202189 239147 217459 239175
rect 217487 239147 217521 239175
rect 217549 239147 232819 239175
rect 232847 239147 232881 239175
rect 232909 239147 248179 239175
rect 248207 239147 248241 239175
rect 248269 239147 263539 239175
rect 263567 239147 263601 239175
rect 263629 239147 278899 239175
rect 278927 239147 278961 239175
rect 278989 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect -958 239113 298990 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 19977 239113
rect 20005 239085 20039 239113
rect 20067 239085 20101 239113
rect 20129 239085 20163 239113
rect 20191 239085 35337 239113
rect 35365 239085 35399 239113
rect 35427 239085 35461 239113
rect 35489 239085 35523 239113
rect 35551 239085 50697 239113
rect 50725 239085 50759 239113
rect 50787 239085 50821 239113
rect 50849 239085 50883 239113
rect 50911 239085 66057 239113
rect 66085 239085 66119 239113
rect 66147 239085 66181 239113
rect 66209 239085 66243 239113
rect 66271 239085 81417 239113
rect 81445 239085 81479 239113
rect 81507 239085 81541 239113
rect 81569 239085 81603 239113
rect 81631 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 109939 239113
rect 109967 239085 110001 239113
rect 110029 239085 125299 239113
rect 125327 239085 125361 239113
rect 125389 239085 140659 239113
rect 140687 239085 140721 239113
rect 140749 239085 156019 239113
rect 156047 239085 156081 239113
rect 156109 239085 171379 239113
rect 171407 239085 171441 239113
rect 171469 239085 186739 239113
rect 186767 239085 186801 239113
rect 186829 239085 202099 239113
rect 202127 239085 202161 239113
rect 202189 239085 217459 239113
rect 217487 239085 217521 239113
rect 217549 239085 232819 239113
rect 232847 239085 232881 239113
rect 232909 239085 248179 239113
rect 248207 239085 248241 239113
rect 248269 239085 263539 239113
rect 263567 239085 263601 239113
rect 263629 239085 278899 239113
rect 278927 239085 278961 239113
rect 278989 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect -958 239051 298990 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 19977 239051
rect 20005 239023 20039 239051
rect 20067 239023 20101 239051
rect 20129 239023 20163 239051
rect 20191 239023 35337 239051
rect 35365 239023 35399 239051
rect 35427 239023 35461 239051
rect 35489 239023 35523 239051
rect 35551 239023 50697 239051
rect 50725 239023 50759 239051
rect 50787 239023 50821 239051
rect 50849 239023 50883 239051
rect 50911 239023 66057 239051
rect 66085 239023 66119 239051
rect 66147 239023 66181 239051
rect 66209 239023 66243 239051
rect 66271 239023 81417 239051
rect 81445 239023 81479 239051
rect 81507 239023 81541 239051
rect 81569 239023 81603 239051
rect 81631 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 109939 239051
rect 109967 239023 110001 239051
rect 110029 239023 125299 239051
rect 125327 239023 125361 239051
rect 125389 239023 140659 239051
rect 140687 239023 140721 239051
rect 140749 239023 156019 239051
rect 156047 239023 156081 239051
rect 156109 239023 171379 239051
rect 171407 239023 171441 239051
rect 171469 239023 186739 239051
rect 186767 239023 186801 239051
rect 186829 239023 202099 239051
rect 202127 239023 202161 239051
rect 202189 239023 217459 239051
rect 217487 239023 217521 239051
rect 217549 239023 232819 239051
rect 232847 239023 232881 239051
rect 232909 239023 248179 239051
rect 248207 239023 248241 239051
rect 248269 239023 263539 239051
rect 263567 239023 263601 239051
rect 263629 239023 278899 239051
rect 278927 239023 278961 239051
rect 278989 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect -958 238989 298990 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 19977 238989
rect 20005 238961 20039 238989
rect 20067 238961 20101 238989
rect 20129 238961 20163 238989
rect 20191 238961 35337 238989
rect 35365 238961 35399 238989
rect 35427 238961 35461 238989
rect 35489 238961 35523 238989
rect 35551 238961 50697 238989
rect 50725 238961 50759 238989
rect 50787 238961 50821 238989
rect 50849 238961 50883 238989
rect 50911 238961 66057 238989
rect 66085 238961 66119 238989
rect 66147 238961 66181 238989
rect 66209 238961 66243 238989
rect 66271 238961 81417 238989
rect 81445 238961 81479 238989
rect 81507 238961 81541 238989
rect 81569 238961 81603 238989
rect 81631 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 109939 238989
rect 109967 238961 110001 238989
rect 110029 238961 125299 238989
rect 125327 238961 125361 238989
rect 125389 238961 140659 238989
rect 140687 238961 140721 238989
rect 140749 238961 156019 238989
rect 156047 238961 156081 238989
rect 156109 238961 171379 238989
rect 171407 238961 171441 238989
rect 171469 238961 186739 238989
rect 186767 238961 186801 238989
rect 186829 238961 202099 238989
rect 202127 238961 202161 238989
rect 202189 238961 217459 238989
rect 217487 238961 217521 238989
rect 217549 238961 232819 238989
rect 232847 238961 232881 238989
rect 232909 238961 248179 238989
rect 248207 238961 248241 238989
rect 248269 238961 263539 238989
rect 263567 238961 263601 238989
rect 263629 238961 278899 238989
rect 278927 238961 278961 238989
rect 278989 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect -958 238913 298990 238961
rect -958 236175 298990 236223
rect -958 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 33477 236175
rect 33505 236147 33539 236175
rect 33567 236147 33601 236175
rect 33629 236147 33663 236175
rect 33691 236147 48837 236175
rect 48865 236147 48899 236175
rect 48927 236147 48961 236175
rect 48989 236147 49023 236175
rect 49051 236147 64197 236175
rect 64225 236147 64259 236175
rect 64287 236147 64321 236175
rect 64349 236147 64383 236175
rect 64411 236147 79557 236175
rect 79585 236147 79619 236175
rect 79647 236147 79681 236175
rect 79709 236147 79743 236175
rect 79771 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 102259 236175
rect 102287 236147 102321 236175
rect 102349 236147 117619 236175
rect 117647 236147 117681 236175
rect 117709 236147 132979 236175
rect 133007 236147 133041 236175
rect 133069 236147 148339 236175
rect 148367 236147 148401 236175
rect 148429 236147 163699 236175
rect 163727 236147 163761 236175
rect 163789 236147 179059 236175
rect 179087 236147 179121 236175
rect 179149 236147 194419 236175
rect 194447 236147 194481 236175
rect 194509 236147 209779 236175
rect 209807 236147 209841 236175
rect 209869 236147 225139 236175
rect 225167 236147 225201 236175
rect 225229 236147 240499 236175
rect 240527 236147 240561 236175
rect 240589 236147 255859 236175
rect 255887 236147 255921 236175
rect 255949 236147 271219 236175
rect 271247 236147 271281 236175
rect 271309 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298990 236175
rect -958 236113 298990 236147
rect -958 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 33477 236113
rect 33505 236085 33539 236113
rect 33567 236085 33601 236113
rect 33629 236085 33663 236113
rect 33691 236085 48837 236113
rect 48865 236085 48899 236113
rect 48927 236085 48961 236113
rect 48989 236085 49023 236113
rect 49051 236085 64197 236113
rect 64225 236085 64259 236113
rect 64287 236085 64321 236113
rect 64349 236085 64383 236113
rect 64411 236085 79557 236113
rect 79585 236085 79619 236113
rect 79647 236085 79681 236113
rect 79709 236085 79743 236113
rect 79771 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 102259 236113
rect 102287 236085 102321 236113
rect 102349 236085 117619 236113
rect 117647 236085 117681 236113
rect 117709 236085 132979 236113
rect 133007 236085 133041 236113
rect 133069 236085 148339 236113
rect 148367 236085 148401 236113
rect 148429 236085 163699 236113
rect 163727 236085 163761 236113
rect 163789 236085 179059 236113
rect 179087 236085 179121 236113
rect 179149 236085 194419 236113
rect 194447 236085 194481 236113
rect 194509 236085 209779 236113
rect 209807 236085 209841 236113
rect 209869 236085 225139 236113
rect 225167 236085 225201 236113
rect 225229 236085 240499 236113
rect 240527 236085 240561 236113
rect 240589 236085 255859 236113
rect 255887 236085 255921 236113
rect 255949 236085 271219 236113
rect 271247 236085 271281 236113
rect 271309 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298990 236113
rect -958 236051 298990 236085
rect -958 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 33477 236051
rect 33505 236023 33539 236051
rect 33567 236023 33601 236051
rect 33629 236023 33663 236051
rect 33691 236023 48837 236051
rect 48865 236023 48899 236051
rect 48927 236023 48961 236051
rect 48989 236023 49023 236051
rect 49051 236023 64197 236051
rect 64225 236023 64259 236051
rect 64287 236023 64321 236051
rect 64349 236023 64383 236051
rect 64411 236023 79557 236051
rect 79585 236023 79619 236051
rect 79647 236023 79681 236051
rect 79709 236023 79743 236051
rect 79771 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 102259 236051
rect 102287 236023 102321 236051
rect 102349 236023 117619 236051
rect 117647 236023 117681 236051
rect 117709 236023 132979 236051
rect 133007 236023 133041 236051
rect 133069 236023 148339 236051
rect 148367 236023 148401 236051
rect 148429 236023 163699 236051
rect 163727 236023 163761 236051
rect 163789 236023 179059 236051
rect 179087 236023 179121 236051
rect 179149 236023 194419 236051
rect 194447 236023 194481 236051
rect 194509 236023 209779 236051
rect 209807 236023 209841 236051
rect 209869 236023 225139 236051
rect 225167 236023 225201 236051
rect 225229 236023 240499 236051
rect 240527 236023 240561 236051
rect 240589 236023 255859 236051
rect 255887 236023 255921 236051
rect 255949 236023 271219 236051
rect 271247 236023 271281 236051
rect 271309 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298990 236051
rect -958 235989 298990 236023
rect -958 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 33477 235989
rect 33505 235961 33539 235989
rect 33567 235961 33601 235989
rect 33629 235961 33663 235989
rect 33691 235961 48837 235989
rect 48865 235961 48899 235989
rect 48927 235961 48961 235989
rect 48989 235961 49023 235989
rect 49051 235961 64197 235989
rect 64225 235961 64259 235989
rect 64287 235961 64321 235989
rect 64349 235961 64383 235989
rect 64411 235961 79557 235989
rect 79585 235961 79619 235989
rect 79647 235961 79681 235989
rect 79709 235961 79743 235989
rect 79771 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 102259 235989
rect 102287 235961 102321 235989
rect 102349 235961 117619 235989
rect 117647 235961 117681 235989
rect 117709 235961 132979 235989
rect 133007 235961 133041 235989
rect 133069 235961 148339 235989
rect 148367 235961 148401 235989
rect 148429 235961 163699 235989
rect 163727 235961 163761 235989
rect 163789 235961 179059 235989
rect 179087 235961 179121 235989
rect 179149 235961 194419 235989
rect 194447 235961 194481 235989
rect 194509 235961 209779 235989
rect 209807 235961 209841 235989
rect 209869 235961 225139 235989
rect 225167 235961 225201 235989
rect 225229 235961 240499 235989
rect 240527 235961 240561 235989
rect 240589 235961 255859 235989
rect 255887 235961 255921 235989
rect 255949 235961 271219 235989
rect 271247 235961 271281 235989
rect 271309 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298990 235989
rect -958 235913 298990 235961
rect -958 230175 298990 230223
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 19977 230175
rect 20005 230147 20039 230175
rect 20067 230147 20101 230175
rect 20129 230147 20163 230175
rect 20191 230147 35337 230175
rect 35365 230147 35399 230175
rect 35427 230147 35461 230175
rect 35489 230147 35523 230175
rect 35551 230147 50697 230175
rect 50725 230147 50759 230175
rect 50787 230147 50821 230175
rect 50849 230147 50883 230175
rect 50911 230147 66057 230175
rect 66085 230147 66119 230175
rect 66147 230147 66181 230175
rect 66209 230147 66243 230175
rect 66271 230147 81417 230175
rect 81445 230147 81479 230175
rect 81507 230147 81541 230175
rect 81569 230147 81603 230175
rect 81631 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 109939 230175
rect 109967 230147 110001 230175
rect 110029 230147 125299 230175
rect 125327 230147 125361 230175
rect 125389 230147 140659 230175
rect 140687 230147 140721 230175
rect 140749 230147 156019 230175
rect 156047 230147 156081 230175
rect 156109 230147 171379 230175
rect 171407 230147 171441 230175
rect 171469 230147 186739 230175
rect 186767 230147 186801 230175
rect 186829 230147 202099 230175
rect 202127 230147 202161 230175
rect 202189 230147 217459 230175
rect 217487 230147 217521 230175
rect 217549 230147 232819 230175
rect 232847 230147 232881 230175
rect 232909 230147 248179 230175
rect 248207 230147 248241 230175
rect 248269 230147 263539 230175
rect 263567 230147 263601 230175
rect 263629 230147 278899 230175
rect 278927 230147 278961 230175
rect 278989 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect -958 230113 298990 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 19977 230113
rect 20005 230085 20039 230113
rect 20067 230085 20101 230113
rect 20129 230085 20163 230113
rect 20191 230085 35337 230113
rect 35365 230085 35399 230113
rect 35427 230085 35461 230113
rect 35489 230085 35523 230113
rect 35551 230085 50697 230113
rect 50725 230085 50759 230113
rect 50787 230085 50821 230113
rect 50849 230085 50883 230113
rect 50911 230085 66057 230113
rect 66085 230085 66119 230113
rect 66147 230085 66181 230113
rect 66209 230085 66243 230113
rect 66271 230085 81417 230113
rect 81445 230085 81479 230113
rect 81507 230085 81541 230113
rect 81569 230085 81603 230113
rect 81631 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 109939 230113
rect 109967 230085 110001 230113
rect 110029 230085 125299 230113
rect 125327 230085 125361 230113
rect 125389 230085 140659 230113
rect 140687 230085 140721 230113
rect 140749 230085 156019 230113
rect 156047 230085 156081 230113
rect 156109 230085 171379 230113
rect 171407 230085 171441 230113
rect 171469 230085 186739 230113
rect 186767 230085 186801 230113
rect 186829 230085 202099 230113
rect 202127 230085 202161 230113
rect 202189 230085 217459 230113
rect 217487 230085 217521 230113
rect 217549 230085 232819 230113
rect 232847 230085 232881 230113
rect 232909 230085 248179 230113
rect 248207 230085 248241 230113
rect 248269 230085 263539 230113
rect 263567 230085 263601 230113
rect 263629 230085 278899 230113
rect 278927 230085 278961 230113
rect 278989 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect -958 230051 298990 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 19977 230051
rect 20005 230023 20039 230051
rect 20067 230023 20101 230051
rect 20129 230023 20163 230051
rect 20191 230023 35337 230051
rect 35365 230023 35399 230051
rect 35427 230023 35461 230051
rect 35489 230023 35523 230051
rect 35551 230023 50697 230051
rect 50725 230023 50759 230051
rect 50787 230023 50821 230051
rect 50849 230023 50883 230051
rect 50911 230023 66057 230051
rect 66085 230023 66119 230051
rect 66147 230023 66181 230051
rect 66209 230023 66243 230051
rect 66271 230023 81417 230051
rect 81445 230023 81479 230051
rect 81507 230023 81541 230051
rect 81569 230023 81603 230051
rect 81631 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 109939 230051
rect 109967 230023 110001 230051
rect 110029 230023 125299 230051
rect 125327 230023 125361 230051
rect 125389 230023 140659 230051
rect 140687 230023 140721 230051
rect 140749 230023 156019 230051
rect 156047 230023 156081 230051
rect 156109 230023 171379 230051
rect 171407 230023 171441 230051
rect 171469 230023 186739 230051
rect 186767 230023 186801 230051
rect 186829 230023 202099 230051
rect 202127 230023 202161 230051
rect 202189 230023 217459 230051
rect 217487 230023 217521 230051
rect 217549 230023 232819 230051
rect 232847 230023 232881 230051
rect 232909 230023 248179 230051
rect 248207 230023 248241 230051
rect 248269 230023 263539 230051
rect 263567 230023 263601 230051
rect 263629 230023 278899 230051
rect 278927 230023 278961 230051
rect 278989 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect -958 229989 298990 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 19977 229989
rect 20005 229961 20039 229989
rect 20067 229961 20101 229989
rect 20129 229961 20163 229989
rect 20191 229961 35337 229989
rect 35365 229961 35399 229989
rect 35427 229961 35461 229989
rect 35489 229961 35523 229989
rect 35551 229961 50697 229989
rect 50725 229961 50759 229989
rect 50787 229961 50821 229989
rect 50849 229961 50883 229989
rect 50911 229961 66057 229989
rect 66085 229961 66119 229989
rect 66147 229961 66181 229989
rect 66209 229961 66243 229989
rect 66271 229961 81417 229989
rect 81445 229961 81479 229989
rect 81507 229961 81541 229989
rect 81569 229961 81603 229989
rect 81631 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 109939 229989
rect 109967 229961 110001 229989
rect 110029 229961 125299 229989
rect 125327 229961 125361 229989
rect 125389 229961 140659 229989
rect 140687 229961 140721 229989
rect 140749 229961 156019 229989
rect 156047 229961 156081 229989
rect 156109 229961 171379 229989
rect 171407 229961 171441 229989
rect 171469 229961 186739 229989
rect 186767 229961 186801 229989
rect 186829 229961 202099 229989
rect 202127 229961 202161 229989
rect 202189 229961 217459 229989
rect 217487 229961 217521 229989
rect 217549 229961 232819 229989
rect 232847 229961 232881 229989
rect 232909 229961 248179 229989
rect 248207 229961 248241 229989
rect 248269 229961 263539 229989
rect 263567 229961 263601 229989
rect 263629 229961 278899 229989
rect 278927 229961 278961 229989
rect 278989 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect -958 229913 298990 229961
rect -958 227175 298990 227223
rect -958 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 33477 227175
rect 33505 227147 33539 227175
rect 33567 227147 33601 227175
rect 33629 227147 33663 227175
rect 33691 227147 48837 227175
rect 48865 227147 48899 227175
rect 48927 227147 48961 227175
rect 48989 227147 49023 227175
rect 49051 227147 64197 227175
rect 64225 227147 64259 227175
rect 64287 227147 64321 227175
rect 64349 227147 64383 227175
rect 64411 227147 79557 227175
rect 79585 227147 79619 227175
rect 79647 227147 79681 227175
rect 79709 227147 79743 227175
rect 79771 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 102259 227175
rect 102287 227147 102321 227175
rect 102349 227147 117619 227175
rect 117647 227147 117681 227175
rect 117709 227147 132979 227175
rect 133007 227147 133041 227175
rect 133069 227147 148339 227175
rect 148367 227147 148401 227175
rect 148429 227147 163699 227175
rect 163727 227147 163761 227175
rect 163789 227147 179059 227175
rect 179087 227147 179121 227175
rect 179149 227147 194419 227175
rect 194447 227147 194481 227175
rect 194509 227147 209779 227175
rect 209807 227147 209841 227175
rect 209869 227147 225139 227175
rect 225167 227147 225201 227175
rect 225229 227147 240499 227175
rect 240527 227147 240561 227175
rect 240589 227147 255859 227175
rect 255887 227147 255921 227175
rect 255949 227147 271219 227175
rect 271247 227147 271281 227175
rect 271309 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298990 227175
rect -958 227113 298990 227147
rect -958 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 33477 227113
rect 33505 227085 33539 227113
rect 33567 227085 33601 227113
rect 33629 227085 33663 227113
rect 33691 227085 48837 227113
rect 48865 227085 48899 227113
rect 48927 227085 48961 227113
rect 48989 227085 49023 227113
rect 49051 227085 64197 227113
rect 64225 227085 64259 227113
rect 64287 227085 64321 227113
rect 64349 227085 64383 227113
rect 64411 227085 79557 227113
rect 79585 227085 79619 227113
rect 79647 227085 79681 227113
rect 79709 227085 79743 227113
rect 79771 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 102259 227113
rect 102287 227085 102321 227113
rect 102349 227085 117619 227113
rect 117647 227085 117681 227113
rect 117709 227085 132979 227113
rect 133007 227085 133041 227113
rect 133069 227085 148339 227113
rect 148367 227085 148401 227113
rect 148429 227085 163699 227113
rect 163727 227085 163761 227113
rect 163789 227085 179059 227113
rect 179087 227085 179121 227113
rect 179149 227085 194419 227113
rect 194447 227085 194481 227113
rect 194509 227085 209779 227113
rect 209807 227085 209841 227113
rect 209869 227085 225139 227113
rect 225167 227085 225201 227113
rect 225229 227085 240499 227113
rect 240527 227085 240561 227113
rect 240589 227085 255859 227113
rect 255887 227085 255921 227113
rect 255949 227085 271219 227113
rect 271247 227085 271281 227113
rect 271309 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298990 227113
rect -958 227051 298990 227085
rect -958 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 33477 227051
rect 33505 227023 33539 227051
rect 33567 227023 33601 227051
rect 33629 227023 33663 227051
rect 33691 227023 48837 227051
rect 48865 227023 48899 227051
rect 48927 227023 48961 227051
rect 48989 227023 49023 227051
rect 49051 227023 64197 227051
rect 64225 227023 64259 227051
rect 64287 227023 64321 227051
rect 64349 227023 64383 227051
rect 64411 227023 79557 227051
rect 79585 227023 79619 227051
rect 79647 227023 79681 227051
rect 79709 227023 79743 227051
rect 79771 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 102259 227051
rect 102287 227023 102321 227051
rect 102349 227023 117619 227051
rect 117647 227023 117681 227051
rect 117709 227023 132979 227051
rect 133007 227023 133041 227051
rect 133069 227023 148339 227051
rect 148367 227023 148401 227051
rect 148429 227023 163699 227051
rect 163727 227023 163761 227051
rect 163789 227023 179059 227051
rect 179087 227023 179121 227051
rect 179149 227023 194419 227051
rect 194447 227023 194481 227051
rect 194509 227023 209779 227051
rect 209807 227023 209841 227051
rect 209869 227023 225139 227051
rect 225167 227023 225201 227051
rect 225229 227023 240499 227051
rect 240527 227023 240561 227051
rect 240589 227023 255859 227051
rect 255887 227023 255921 227051
rect 255949 227023 271219 227051
rect 271247 227023 271281 227051
rect 271309 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298990 227051
rect -958 226989 298990 227023
rect -958 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 33477 226989
rect 33505 226961 33539 226989
rect 33567 226961 33601 226989
rect 33629 226961 33663 226989
rect 33691 226961 48837 226989
rect 48865 226961 48899 226989
rect 48927 226961 48961 226989
rect 48989 226961 49023 226989
rect 49051 226961 64197 226989
rect 64225 226961 64259 226989
rect 64287 226961 64321 226989
rect 64349 226961 64383 226989
rect 64411 226961 79557 226989
rect 79585 226961 79619 226989
rect 79647 226961 79681 226989
rect 79709 226961 79743 226989
rect 79771 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 102259 226989
rect 102287 226961 102321 226989
rect 102349 226961 117619 226989
rect 117647 226961 117681 226989
rect 117709 226961 132979 226989
rect 133007 226961 133041 226989
rect 133069 226961 148339 226989
rect 148367 226961 148401 226989
rect 148429 226961 163699 226989
rect 163727 226961 163761 226989
rect 163789 226961 179059 226989
rect 179087 226961 179121 226989
rect 179149 226961 194419 226989
rect 194447 226961 194481 226989
rect 194509 226961 209779 226989
rect 209807 226961 209841 226989
rect 209869 226961 225139 226989
rect 225167 226961 225201 226989
rect 225229 226961 240499 226989
rect 240527 226961 240561 226989
rect 240589 226961 255859 226989
rect 255887 226961 255921 226989
rect 255949 226961 271219 226989
rect 271247 226961 271281 226989
rect 271309 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298990 226989
rect -958 226913 298990 226961
rect -958 221175 298990 221223
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 19977 221175
rect 20005 221147 20039 221175
rect 20067 221147 20101 221175
rect 20129 221147 20163 221175
rect 20191 221147 35337 221175
rect 35365 221147 35399 221175
rect 35427 221147 35461 221175
rect 35489 221147 35523 221175
rect 35551 221147 50697 221175
rect 50725 221147 50759 221175
rect 50787 221147 50821 221175
rect 50849 221147 50883 221175
rect 50911 221147 66057 221175
rect 66085 221147 66119 221175
rect 66147 221147 66181 221175
rect 66209 221147 66243 221175
rect 66271 221147 81417 221175
rect 81445 221147 81479 221175
rect 81507 221147 81541 221175
rect 81569 221147 81603 221175
rect 81631 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 109939 221175
rect 109967 221147 110001 221175
rect 110029 221147 125299 221175
rect 125327 221147 125361 221175
rect 125389 221147 140659 221175
rect 140687 221147 140721 221175
rect 140749 221147 156019 221175
rect 156047 221147 156081 221175
rect 156109 221147 171379 221175
rect 171407 221147 171441 221175
rect 171469 221147 186739 221175
rect 186767 221147 186801 221175
rect 186829 221147 202099 221175
rect 202127 221147 202161 221175
rect 202189 221147 217459 221175
rect 217487 221147 217521 221175
rect 217549 221147 232819 221175
rect 232847 221147 232881 221175
rect 232909 221147 248179 221175
rect 248207 221147 248241 221175
rect 248269 221147 263539 221175
rect 263567 221147 263601 221175
rect 263629 221147 278899 221175
rect 278927 221147 278961 221175
rect 278989 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect -958 221113 298990 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 19977 221113
rect 20005 221085 20039 221113
rect 20067 221085 20101 221113
rect 20129 221085 20163 221113
rect 20191 221085 35337 221113
rect 35365 221085 35399 221113
rect 35427 221085 35461 221113
rect 35489 221085 35523 221113
rect 35551 221085 50697 221113
rect 50725 221085 50759 221113
rect 50787 221085 50821 221113
rect 50849 221085 50883 221113
rect 50911 221085 66057 221113
rect 66085 221085 66119 221113
rect 66147 221085 66181 221113
rect 66209 221085 66243 221113
rect 66271 221085 81417 221113
rect 81445 221085 81479 221113
rect 81507 221085 81541 221113
rect 81569 221085 81603 221113
rect 81631 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 109939 221113
rect 109967 221085 110001 221113
rect 110029 221085 125299 221113
rect 125327 221085 125361 221113
rect 125389 221085 140659 221113
rect 140687 221085 140721 221113
rect 140749 221085 156019 221113
rect 156047 221085 156081 221113
rect 156109 221085 171379 221113
rect 171407 221085 171441 221113
rect 171469 221085 186739 221113
rect 186767 221085 186801 221113
rect 186829 221085 202099 221113
rect 202127 221085 202161 221113
rect 202189 221085 217459 221113
rect 217487 221085 217521 221113
rect 217549 221085 232819 221113
rect 232847 221085 232881 221113
rect 232909 221085 248179 221113
rect 248207 221085 248241 221113
rect 248269 221085 263539 221113
rect 263567 221085 263601 221113
rect 263629 221085 278899 221113
rect 278927 221085 278961 221113
rect 278989 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect -958 221051 298990 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 19977 221051
rect 20005 221023 20039 221051
rect 20067 221023 20101 221051
rect 20129 221023 20163 221051
rect 20191 221023 35337 221051
rect 35365 221023 35399 221051
rect 35427 221023 35461 221051
rect 35489 221023 35523 221051
rect 35551 221023 50697 221051
rect 50725 221023 50759 221051
rect 50787 221023 50821 221051
rect 50849 221023 50883 221051
rect 50911 221023 66057 221051
rect 66085 221023 66119 221051
rect 66147 221023 66181 221051
rect 66209 221023 66243 221051
rect 66271 221023 81417 221051
rect 81445 221023 81479 221051
rect 81507 221023 81541 221051
rect 81569 221023 81603 221051
rect 81631 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 109939 221051
rect 109967 221023 110001 221051
rect 110029 221023 125299 221051
rect 125327 221023 125361 221051
rect 125389 221023 140659 221051
rect 140687 221023 140721 221051
rect 140749 221023 156019 221051
rect 156047 221023 156081 221051
rect 156109 221023 171379 221051
rect 171407 221023 171441 221051
rect 171469 221023 186739 221051
rect 186767 221023 186801 221051
rect 186829 221023 202099 221051
rect 202127 221023 202161 221051
rect 202189 221023 217459 221051
rect 217487 221023 217521 221051
rect 217549 221023 232819 221051
rect 232847 221023 232881 221051
rect 232909 221023 248179 221051
rect 248207 221023 248241 221051
rect 248269 221023 263539 221051
rect 263567 221023 263601 221051
rect 263629 221023 278899 221051
rect 278927 221023 278961 221051
rect 278989 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect -958 220989 298990 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 19977 220989
rect 20005 220961 20039 220989
rect 20067 220961 20101 220989
rect 20129 220961 20163 220989
rect 20191 220961 35337 220989
rect 35365 220961 35399 220989
rect 35427 220961 35461 220989
rect 35489 220961 35523 220989
rect 35551 220961 50697 220989
rect 50725 220961 50759 220989
rect 50787 220961 50821 220989
rect 50849 220961 50883 220989
rect 50911 220961 66057 220989
rect 66085 220961 66119 220989
rect 66147 220961 66181 220989
rect 66209 220961 66243 220989
rect 66271 220961 81417 220989
rect 81445 220961 81479 220989
rect 81507 220961 81541 220989
rect 81569 220961 81603 220989
rect 81631 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 109939 220989
rect 109967 220961 110001 220989
rect 110029 220961 125299 220989
rect 125327 220961 125361 220989
rect 125389 220961 140659 220989
rect 140687 220961 140721 220989
rect 140749 220961 156019 220989
rect 156047 220961 156081 220989
rect 156109 220961 171379 220989
rect 171407 220961 171441 220989
rect 171469 220961 186739 220989
rect 186767 220961 186801 220989
rect 186829 220961 202099 220989
rect 202127 220961 202161 220989
rect 202189 220961 217459 220989
rect 217487 220961 217521 220989
rect 217549 220961 232819 220989
rect 232847 220961 232881 220989
rect 232909 220961 248179 220989
rect 248207 220961 248241 220989
rect 248269 220961 263539 220989
rect 263567 220961 263601 220989
rect 263629 220961 278899 220989
rect 278927 220961 278961 220989
rect 278989 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect -958 220913 298990 220961
rect -958 218175 298990 218223
rect -958 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 33477 218175
rect 33505 218147 33539 218175
rect 33567 218147 33601 218175
rect 33629 218147 33663 218175
rect 33691 218147 48837 218175
rect 48865 218147 48899 218175
rect 48927 218147 48961 218175
rect 48989 218147 49023 218175
rect 49051 218147 64197 218175
rect 64225 218147 64259 218175
rect 64287 218147 64321 218175
rect 64349 218147 64383 218175
rect 64411 218147 79557 218175
rect 79585 218147 79619 218175
rect 79647 218147 79681 218175
rect 79709 218147 79743 218175
rect 79771 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 102259 218175
rect 102287 218147 102321 218175
rect 102349 218147 117619 218175
rect 117647 218147 117681 218175
rect 117709 218147 132979 218175
rect 133007 218147 133041 218175
rect 133069 218147 148339 218175
rect 148367 218147 148401 218175
rect 148429 218147 163699 218175
rect 163727 218147 163761 218175
rect 163789 218147 179059 218175
rect 179087 218147 179121 218175
rect 179149 218147 194419 218175
rect 194447 218147 194481 218175
rect 194509 218147 209779 218175
rect 209807 218147 209841 218175
rect 209869 218147 225139 218175
rect 225167 218147 225201 218175
rect 225229 218147 240499 218175
rect 240527 218147 240561 218175
rect 240589 218147 255859 218175
rect 255887 218147 255921 218175
rect 255949 218147 271219 218175
rect 271247 218147 271281 218175
rect 271309 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298990 218175
rect -958 218113 298990 218147
rect -958 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 33477 218113
rect 33505 218085 33539 218113
rect 33567 218085 33601 218113
rect 33629 218085 33663 218113
rect 33691 218085 48837 218113
rect 48865 218085 48899 218113
rect 48927 218085 48961 218113
rect 48989 218085 49023 218113
rect 49051 218085 64197 218113
rect 64225 218085 64259 218113
rect 64287 218085 64321 218113
rect 64349 218085 64383 218113
rect 64411 218085 79557 218113
rect 79585 218085 79619 218113
rect 79647 218085 79681 218113
rect 79709 218085 79743 218113
rect 79771 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 102259 218113
rect 102287 218085 102321 218113
rect 102349 218085 117619 218113
rect 117647 218085 117681 218113
rect 117709 218085 132979 218113
rect 133007 218085 133041 218113
rect 133069 218085 148339 218113
rect 148367 218085 148401 218113
rect 148429 218085 163699 218113
rect 163727 218085 163761 218113
rect 163789 218085 179059 218113
rect 179087 218085 179121 218113
rect 179149 218085 194419 218113
rect 194447 218085 194481 218113
rect 194509 218085 209779 218113
rect 209807 218085 209841 218113
rect 209869 218085 225139 218113
rect 225167 218085 225201 218113
rect 225229 218085 240499 218113
rect 240527 218085 240561 218113
rect 240589 218085 255859 218113
rect 255887 218085 255921 218113
rect 255949 218085 271219 218113
rect 271247 218085 271281 218113
rect 271309 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298990 218113
rect -958 218051 298990 218085
rect -958 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 33477 218051
rect 33505 218023 33539 218051
rect 33567 218023 33601 218051
rect 33629 218023 33663 218051
rect 33691 218023 48837 218051
rect 48865 218023 48899 218051
rect 48927 218023 48961 218051
rect 48989 218023 49023 218051
rect 49051 218023 64197 218051
rect 64225 218023 64259 218051
rect 64287 218023 64321 218051
rect 64349 218023 64383 218051
rect 64411 218023 79557 218051
rect 79585 218023 79619 218051
rect 79647 218023 79681 218051
rect 79709 218023 79743 218051
rect 79771 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 102259 218051
rect 102287 218023 102321 218051
rect 102349 218023 117619 218051
rect 117647 218023 117681 218051
rect 117709 218023 132979 218051
rect 133007 218023 133041 218051
rect 133069 218023 148339 218051
rect 148367 218023 148401 218051
rect 148429 218023 163699 218051
rect 163727 218023 163761 218051
rect 163789 218023 179059 218051
rect 179087 218023 179121 218051
rect 179149 218023 194419 218051
rect 194447 218023 194481 218051
rect 194509 218023 209779 218051
rect 209807 218023 209841 218051
rect 209869 218023 225139 218051
rect 225167 218023 225201 218051
rect 225229 218023 240499 218051
rect 240527 218023 240561 218051
rect 240589 218023 255859 218051
rect 255887 218023 255921 218051
rect 255949 218023 271219 218051
rect 271247 218023 271281 218051
rect 271309 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298990 218051
rect -958 217989 298990 218023
rect -958 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 33477 217989
rect 33505 217961 33539 217989
rect 33567 217961 33601 217989
rect 33629 217961 33663 217989
rect 33691 217961 48837 217989
rect 48865 217961 48899 217989
rect 48927 217961 48961 217989
rect 48989 217961 49023 217989
rect 49051 217961 64197 217989
rect 64225 217961 64259 217989
rect 64287 217961 64321 217989
rect 64349 217961 64383 217989
rect 64411 217961 79557 217989
rect 79585 217961 79619 217989
rect 79647 217961 79681 217989
rect 79709 217961 79743 217989
rect 79771 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 102259 217989
rect 102287 217961 102321 217989
rect 102349 217961 117619 217989
rect 117647 217961 117681 217989
rect 117709 217961 132979 217989
rect 133007 217961 133041 217989
rect 133069 217961 148339 217989
rect 148367 217961 148401 217989
rect 148429 217961 163699 217989
rect 163727 217961 163761 217989
rect 163789 217961 179059 217989
rect 179087 217961 179121 217989
rect 179149 217961 194419 217989
rect 194447 217961 194481 217989
rect 194509 217961 209779 217989
rect 209807 217961 209841 217989
rect 209869 217961 225139 217989
rect 225167 217961 225201 217989
rect 225229 217961 240499 217989
rect 240527 217961 240561 217989
rect 240589 217961 255859 217989
rect 255887 217961 255921 217989
rect 255949 217961 271219 217989
rect 271247 217961 271281 217989
rect 271309 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298990 217989
rect -958 217913 298990 217961
rect -958 212175 298990 212223
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 19977 212175
rect 20005 212147 20039 212175
rect 20067 212147 20101 212175
rect 20129 212147 20163 212175
rect 20191 212147 35337 212175
rect 35365 212147 35399 212175
rect 35427 212147 35461 212175
rect 35489 212147 35523 212175
rect 35551 212147 50697 212175
rect 50725 212147 50759 212175
rect 50787 212147 50821 212175
rect 50849 212147 50883 212175
rect 50911 212147 66057 212175
rect 66085 212147 66119 212175
rect 66147 212147 66181 212175
rect 66209 212147 66243 212175
rect 66271 212147 81417 212175
rect 81445 212147 81479 212175
rect 81507 212147 81541 212175
rect 81569 212147 81603 212175
rect 81631 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 109939 212175
rect 109967 212147 110001 212175
rect 110029 212147 125299 212175
rect 125327 212147 125361 212175
rect 125389 212147 140659 212175
rect 140687 212147 140721 212175
rect 140749 212147 156019 212175
rect 156047 212147 156081 212175
rect 156109 212147 171379 212175
rect 171407 212147 171441 212175
rect 171469 212147 186739 212175
rect 186767 212147 186801 212175
rect 186829 212147 202099 212175
rect 202127 212147 202161 212175
rect 202189 212147 217459 212175
rect 217487 212147 217521 212175
rect 217549 212147 232819 212175
rect 232847 212147 232881 212175
rect 232909 212147 248179 212175
rect 248207 212147 248241 212175
rect 248269 212147 263539 212175
rect 263567 212147 263601 212175
rect 263629 212147 278899 212175
rect 278927 212147 278961 212175
rect 278989 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect -958 212113 298990 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 19977 212113
rect 20005 212085 20039 212113
rect 20067 212085 20101 212113
rect 20129 212085 20163 212113
rect 20191 212085 35337 212113
rect 35365 212085 35399 212113
rect 35427 212085 35461 212113
rect 35489 212085 35523 212113
rect 35551 212085 50697 212113
rect 50725 212085 50759 212113
rect 50787 212085 50821 212113
rect 50849 212085 50883 212113
rect 50911 212085 66057 212113
rect 66085 212085 66119 212113
rect 66147 212085 66181 212113
rect 66209 212085 66243 212113
rect 66271 212085 81417 212113
rect 81445 212085 81479 212113
rect 81507 212085 81541 212113
rect 81569 212085 81603 212113
rect 81631 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 109939 212113
rect 109967 212085 110001 212113
rect 110029 212085 125299 212113
rect 125327 212085 125361 212113
rect 125389 212085 140659 212113
rect 140687 212085 140721 212113
rect 140749 212085 156019 212113
rect 156047 212085 156081 212113
rect 156109 212085 171379 212113
rect 171407 212085 171441 212113
rect 171469 212085 186739 212113
rect 186767 212085 186801 212113
rect 186829 212085 202099 212113
rect 202127 212085 202161 212113
rect 202189 212085 217459 212113
rect 217487 212085 217521 212113
rect 217549 212085 232819 212113
rect 232847 212085 232881 212113
rect 232909 212085 248179 212113
rect 248207 212085 248241 212113
rect 248269 212085 263539 212113
rect 263567 212085 263601 212113
rect 263629 212085 278899 212113
rect 278927 212085 278961 212113
rect 278989 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect -958 212051 298990 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 19977 212051
rect 20005 212023 20039 212051
rect 20067 212023 20101 212051
rect 20129 212023 20163 212051
rect 20191 212023 35337 212051
rect 35365 212023 35399 212051
rect 35427 212023 35461 212051
rect 35489 212023 35523 212051
rect 35551 212023 50697 212051
rect 50725 212023 50759 212051
rect 50787 212023 50821 212051
rect 50849 212023 50883 212051
rect 50911 212023 66057 212051
rect 66085 212023 66119 212051
rect 66147 212023 66181 212051
rect 66209 212023 66243 212051
rect 66271 212023 81417 212051
rect 81445 212023 81479 212051
rect 81507 212023 81541 212051
rect 81569 212023 81603 212051
rect 81631 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 109939 212051
rect 109967 212023 110001 212051
rect 110029 212023 125299 212051
rect 125327 212023 125361 212051
rect 125389 212023 140659 212051
rect 140687 212023 140721 212051
rect 140749 212023 156019 212051
rect 156047 212023 156081 212051
rect 156109 212023 171379 212051
rect 171407 212023 171441 212051
rect 171469 212023 186739 212051
rect 186767 212023 186801 212051
rect 186829 212023 202099 212051
rect 202127 212023 202161 212051
rect 202189 212023 217459 212051
rect 217487 212023 217521 212051
rect 217549 212023 232819 212051
rect 232847 212023 232881 212051
rect 232909 212023 248179 212051
rect 248207 212023 248241 212051
rect 248269 212023 263539 212051
rect 263567 212023 263601 212051
rect 263629 212023 278899 212051
rect 278927 212023 278961 212051
rect 278989 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect -958 211989 298990 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 19977 211989
rect 20005 211961 20039 211989
rect 20067 211961 20101 211989
rect 20129 211961 20163 211989
rect 20191 211961 35337 211989
rect 35365 211961 35399 211989
rect 35427 211961 35461 211989
rect 35489 211961 35523 211989
rect 35551 211961 50697 211989
rect 50725 211961 50759 211989
rect 50787 211961 50821 211989
rect 50849 211961 50883 211989
rect 50911 211961 66057 211989
rect 66085 211961 66119 211989
rect 66147 211961 66181 211989
rect 66209 211961 66243 211989
rect 66271 211961 81417 211989
rect 81445 211961 81479 211989
rect 81507 211961 81541 211989
rect 81569 211961 81603 211989
rect 81631 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 109939 211989
rect 109967 211961 110001 211989
rect 110029 211961 125299 211989
rect 125327 211961 125361 211989
rect 125389 211961 140659 211989
rect 140687 211961 140721 211989
rect 140749 211961 156019 211989
rect 156047 211961 156081 211989
rect 156109 211961 171379 211989
rect 171407 211961 171441 211989
rect 171469 211961 186739 211989
rect 186767 211961 186801 211989
rect 186829 211961 202099 211989
rect 202127 211961 202161 211989
rect 202189 211961 217459 211989
rect 217487 211961 217521 211989
rect 217549 211961 232819 211989
rect 232847 211961 232881 211989
rect 232909 211961 248179 211989
rect 248207 211961 248241 211989
rect 248269 211961 263539 211989
rect 263567 211961 263601 211989
rect 263629 211961 278899 211989
rect 278927 211961 278961 211989
rect 278989 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect -958 211913 298990 211961
rect -958 209175 298990 209223
rect -958 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 33477 209175
rect 33505 209147 33539 209175
rect 33567 209147 33601 209175
rect 33629 209147 33663 209175
rect 33691 209147 48837 209175
rect 48865 209147 48899 209175
rect 48927 209147 48961 209175
rect 48989 209147 49023 209175
rect 49051 209147 64197 209175
rect 64225 209147 64259 209175
rect 64287 209147 64321 209175
rect 64349 209147 64383 209175
rect 64411 209147 79557 209175
rect 79585 209147 79619 209175
rect 79647 209147 79681 209175
rect 79709 209147 79743 209175
rect 79771 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 102259 209175
rect 102287 209147 102321 209175
rect 102349 209147 117619 209175
rect 117647 209147 117681 209175
rect 117709 209147 132979 209175
rect 133007 209147 133041 209175
rect 133069 209147 148339 209175
rect 148367 209147 148401 209175
rect 148429 209147 163699 209175
rect 163727 209147 163761 209175
rect 163789 209147 179059 209175
rect 179087 209147 179121 209175
rect 179149 209147 194419 209175
rect 194447 209147 194481 209175
rect 194509 209147 209779 209175
rect 209807 209147 209841 209175
rect 209869 209147 225139 209175
rect 225167 209147 225201 209175
rect 225229 209147 240499 209175
rect 240527 209147 240561 209175
rect 240589 209147 255859 209175
rect 255887 209147 255921 209175
rect 255949 209147 271219 209175
rect 271247 209147 271281 209175
rect 271309 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298990 209175
rect -958 209113 298990 209147
rect -958 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 33477 209113
rect 33505 209085 33539 209113
rect 33567 209085 33601 209113
rect 33629 209085 33663 209113
rect 33691 209085 48837 209113
rect 48865 209085 48899 209113
rect 48927 209085 48961 209113
rect 48989 209085 49023 209113
rect 49051 209085 64197 209113
rect 64225 209085 64259 209113
rect 64287 209085 64321 209113
rect 64349 209085 64383 209113
rect 64411 209085 79557 209113
rect 79585 209085 79619 209113
rect 79647 209085 79681 209113
rect 79709 209085 79743 209113
rect 79771 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 102259 209113
rect 102287 209085 102321 209113
rect 102349 209085 117619 209113
rect 117647 209085 117681 209113
rect 117709 209085 132979 209113
rect 133007 209085 133041 209113
rect 133069 209085 148339 209113
rect 148367 209085 148401 209113
rect 148429 209085 163699 209113
rect 163727 209085 163761 209113
rect 163789 209085 179059 209113
rect 179087 209085 179121 209113
rect 179149 209085 194419 209113
rect 194447 209085 194481 209113
rect 194509 209085 209779 209113
rect 209807 209085 209841 209113
rect 209869 209085 225139 209113
rect 225167 209085 225201 209113
rect 225229 209085 240499 209113
rect 240527 209085 240561 209113
rect 240589 209085 255859 209113
rect 255887 209085 255921 209113
rect 255949 209085 271219 209113
rect 271247 209085 271281 209113
rect 271309 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298990 209113
rect -958 209051 298990 209085
rect -958 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 33477 209051
rect 33505 209023 33539 209051
rect 33567 209023 33601 209051
rect 33629 209023 33663 209051
rect 33691 209023 48837 209051
rect 48865 209023 48899 209051
rect 48927 209023 48961 209051
rect 48989 209023 49023 209051
rect 49051 209023 64197 209051
rect 64225 209023 64259 209051
rect 64287 209023 64321 209051
rect 64349 209023 64383 209051
rect 64411 209023 79557 209051
rect 79585 209023 79619 209051
rect 79647 209023 79681 209051
rect 79709 209023 79743 209051
rect 79771 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 102259 209051
rect 102287 209023 102321 209051
rect 102349 209023 117619 209051
rect 117647 209023 117681 209051
rect 117709 209023 132979 209051
rect 133007 209023 133041 209051
rect 133069 209023 148339 209051
rect 148367 209023 148401 209051
rect 148429 209023 163699 209051
rect 163727 209023 163761 209051
rect 163789 209023 179059 209051
rect 179087 209023 179121 209051
rect 179149 209023 194419 209051
rect 194447 209023 194481 209051
rect 194509 209023 209779 209051
rect 209807 209023 209841 209051
rect 209869 209023 225139 209051
rect 225167 209023 225201 209051
rect 225229 209023 240499 209051
rect 240527 209023 240561 209051
rect 240589 209023 255859 209051
rect 255887 209023 255921 209051
rect 255949 209023 271219 209051
rect 271247 209023 271281 209051
rect 271309 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298990 209051
rect -958 208989 298990 209023
rect -958 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 33477 208989
rect 33505 208961 33539 208989
rect 33567 208961 33601 208989
rect 33629 208961 33663 208989
rect 33691 208961 48837 208989
rect 48865 208961 48899 208989
rect 48927 208961 48961 208989
rect 48989 208961 49023 208989
rect 49051 208961 64197 208989
rect 64225 208961 64259 208989
rect 64287 208961 64321 208989
rect 64349 208961 64383 208989
rect 64411 208961 79557 208989
rect 79585 208961 79619 208989
rect 79647 208961 79681 208989
rect 79709 208961 79743 208989
rect 79771 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 102259 208989
rect 102287 208961 102321 208989
rect 102349 208961 117619 208989
rect 117647 208961 117681 208989
rect 117709 208961 132979 208989
rect 133007 208961 133041 208989
rect 133069 208961 148339 208989
rect 148367 208961 148401 208989
rect 148429 208961 163699 208989
rect 163727 208961 163761 208989
rect 163789 208961 179059 208989
rect 179087 208961 179121 208989
rect 179149 208961 194419 208989
rect 194447 208961 194481 208989
rect 194509 208961 209779 208989
rect 209807 208961 209841 208989
rect 209869 208961 225139 208989
rect 225167 208961 225201 208989
rect 225229 208961 240499 208989
rect 240527 208961 240561 208989
rect 240589 208961 255859 208989
rect 255887 208961 255921 208989
rect 255949 208961 271219 208989
rect 271247 208961 271281 208989
rect 271309 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298990 208989
rect -958 208913 298990 208961
rect -958 203175 298990 203223
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 19977 203175
rect 20005 203147 20039 203175
rect 20067 203147 20101 203175
rect 20129 203147 20163 203175
rect 20191 203147 35337 203175
rect 35365 203147 35399 203175
rect 35427 203147 35461 203175
rect 35489 203147 35523 203175
rect 35551 203147 50697 203175
rect 50725 203147 50759 203175
rect 50787 203147 50821 203175
rect 50849 203147 50883 203175
rect 50911 203147 66057 203175
rect 66085 203147 66119 203175
rect 66147 203147 66181 203175
rect 66209 203147 66243 203175
rect 66271 203147 81417 203175
rect 81445 203147 81479 203175
rect 81507 203147 81541 203175
rect 81569 203147 81603 203175
rect 81631 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 109939 203175
rect 109967 203147 110001 203175
rect 110029 203147 125299 203175
rect 125327 203147 125361 203175
rect 125389 203147 140659 203175
rect 140687 203147 140721 203175
rect 140749 203147 156019 203175
rect 156047 203147 156081 203175
rect 156109 203147 171379 203175
rect 171407 203147 171441 203175
rect 171469 203147 186739 203175
rect 186767 203147 186801 203175
rect 186829 203147 202099 203175
rect 202127 203147 202161 203175
rect 202189 203147 217459 203175
rect 217487 203147 217521 203175
rect 217549 203147 232819 203175
rect 232847 203147 232881 203175
rect 232909 203147 248179 203175
rect 248207 203147 248241 203175
rect 248269 203147 263539 203175
rect 263567 203147 263601 203175
rect 263629 203147 278899 203175
rect 278927 203147 278961 203175
rect 278989 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect -958 203113 298990 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 19977 203113
rect 20005 203085 20039 203113
rect 20067 203085 20101 203113
rect 20129 203085 20163 203113
rect 20191 203085 35337 203113
rect 35365 203085 35399 203113
rect 35427 203085 35461 203113
rect 35489 203085 35523 203113
rect 35551 203085 50697 203113
rect 50725 203085 50759 203113
rect 50787 203085 50821 203113
rect 50849 203085 50883 203113
rect 50911 203085 66057 203113
rect 66085 203085 66119 203113
rect 66147 203085 66181 203113
rect 66209 203085 66243 203113
rect 66271 203085 81417 203113
rect 81445 203085 81479 203113
rect 81507 203085 81541 203113
rect 81569 203085 81603 203113
rect 81631 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 109939 203113
rect 109967 203085 110001 203113
rect 110029 203085 125299 203113
rect 125327 203085 125361 203113
rect 125389 203085 140659 203113
rect 140687 203085 140721 203113
rect 140749 203085 156019 203113
rect 156047 203085 156081 203113
rect 156109 203085 171379 203113
rect 171407 203085 171441 203113
rect 171469 203085 186739 203113
rect 186767 203085 186801 203113
rect 186829 203085 202099 203113
rect 202127 203085 202161 203113
rect 202189 203085 217459 203113
rect 217487 203085 217521 203113
rect 217549 203085 232819 203113
rect 232847 203085 232881 203113
rect 232909 203085 248179 203113
rect 248207 203085 248241 203113
rect 248269 203085 263539 203113
rect 263567 203085 263601 203113
rect 263629 203085 278899 203113
rect 278927 203085 278961 203113
rect 278989 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect -958 203051 298990 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 19977 203051
rect 20005 203023 20039 203051
rect 20067 203023 20101 203051
rect 20129 203023 20163 203051
rect 20191 203023 35337 203051
rect 35365 203023 35399 203051
rect 35427 203023 35461 203051
rect 35489 203023 35523 203051
rect 35551 203023 50697 203051
rect 50725 203023 50759 203051
rect 50787 203023 50821 203051
rect 50849 203023 50883 203051
rect 50911 203023 66057 203051
rect 66085 203023 66119 203051
rect 66147 203023 66181 203051
rect 66209 203023 66243 203051
rect 66271 203023 81417 203051
rect 81445 203023 81479 203051
rect 81507 203023 81541 203051
rect 81569 203023 81603 203051
rect 81631 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 109939 203051
rect 109967 203023 110001 203051
rect 110029 203023 125299 203051
rect 125327 203023 125361 203051
rect 125389 203023 140659 203051
rect 140687 203023 140721 203051
rect 140749 203023 156019 203051
rect 156047 203023 156081 203051
rect 156109 203023 171379 203051
rect 171407 203023 171441 203051
rect 171469 203023 186739 203051
rect 186767 203023 186801 203051
rect 186829 203023 202099 203051
rect 202127 203023 202161 203051
rect 202189 203023 217459 203051
rect 217487 203023 217521 203051
rect 217549 203023 232819 203051
rect 232847 203023 232881 203051
rect 232909 203023 248179 203051
rect 248207 203023 248241 203051
rect 248269 203023 263539 203051
rect 263567 203023 263601 203051
rect 263629 203023 278899 203051
rect 278927 203023 278961 203051
rect 278989 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect -958 202989 298990 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 19977 202989
rect 20005 202961 20039 202989
rect 20067 202961 20101 202989
rect 20129 202961 20163 202989
rect 20191 202961 35337 202989
rect 35365 202961 35399 202989
rect 35427 202961 35461 202989
rect 35489 202961 35523 202989
rect 35551 202961 50697 202989
rect 50725 202961 50759 202989
rect 50787 202961 50821 202989
rect 50849 202961 50883 202989
rect 50911 202961 66057 202989
rect 66085 202961 66119 202989
rect 66147 202961 66181 202989
rect 66209 202961 66243 202989
rect 66271 202961 81417 202989
rect 81445 202961 81479 202989
rect 81507 202961 81541 202989
rect 81569 202961 81603 202989
rect 81631 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 109939 202989
rect 109967 202961 110001 202989
rect 110029 202961 125299 202989
rect 125327 202961 125361 202989
rect 125389 202961 140659 202989
rect 140687 202961 140721 202989
rect 140749 202961 156019 202989
rect 156047 202961 156081 202989
rect 156109 202961 171379 202989
rect 171407 202961 171441 202989
rect 171469 202961 186739 202989
rect 186767 202961 186801 202989
rect 186829 202961 202099 202989
rect 202127 202961 202161 202989
rect 202189 202961 217459 202989
rect 217487 202961 217521 202989
rect 217549 202961 232819 202989
rect 232847 202961 232881 202989
rect 232909 202961 248179 202989
rect 248207 202961 248241 202989
rect 248269 202961 263539 202989
rect 263567 202961 263601 202989
rect 263629 202961 278899 202989
rect 278927 202961 278961 202989
rect 278989 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect -958 202913 298990 202961
rect -958 200175 298990 200223
rect -958 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 33477 200175
rect 33505 200147 33539 200175
rect 33567 200147 33601 200175
rect 33629 200147 33663 200175
rect 33691 200147 48837 200175
rect 48865 200147 48899 200175
rect 48927 200147 48961 200175
rect 48989 200147 49023 200175
rect 49051 200147 64197 200175
rect 64225 200147 64259 200175
rect 64287 200147 64321 200175
rect 64349 200147 64383 200175
rect 64411 200147 79557 200175
rect 79585 200147 79619 200175
rect 79647 200147 79681 200175
rect 79709 200147 79743 200175
rect 79771 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 102259 200175
rect 102287 200147 102321 200175
rect 102349 200147 117619 200175
rect 117647 200147 117681 200175
rect 117709 200147 132979 200175
rect 133007 200147 133041 200175
rect 133069 200147 148339 200175
rect 148367 200147 148401 200175
rect 148429 200147 163699 200175
rect 163727 200147 163761 200175
rect 163789 200147 179059 200175
rect 179087 200147 179121 200175
rect 179149 200147 194419 200175
rect 194447 200147 194481 200175
rect 194509 200147 209779 200175
rect 209807 200147 209841 200175
rect 209869 200147 225139 200175
rect 225167 200147 225201 200175
rect 225229 200147 240499 200175
rect 240527 200147 240561 200175
rect 240589 200147 255859 200175
rect 255887 200147 255921 200175
rect 255949 200147 271219 200175
rect 271247 200147 271281 200175
rect 271309 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298990 200175
rect -958 200113 298990 200147
rect -958 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 33477 200113
rect 33505 200085 33539 200113
rect 33567 200085 33601 200113
rect 33629 200085 33663 200113
rect 33691 200085 48837 200113
rect 48865 200085 48899 200113
rect 48927 200085 48961 200113
rect 48989 200085 49023 200113
rect 49051 200085 64197 200113
rect 64225 200085 64259 200113
rect 64287 200085 64321 200113
rect 64349 200085 64383 200113
rect 64411 200085 79557 200113
rect 79585 200085 79619 200113
rect 79647 200085 79681 200113
rect 79709 200085 79743 200113
rect 79771 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 102259 200113
rect 102287 200085 102321 200113
rect 102349 200085 117619 200113
rect 117647 200085 117681 200113
rect 117709 200085 132979 200113
rect 133007 200085 133041 200113
rect 133069 200085 148339 200113
rect 148367 200085 148401 200113
rect 148429 200085 163699 200113
rect 163727 200085 163761 200113
rect 163789 200085 179059 200113
rect 179087 200085 179121 200113
rect 179149 200085 194419 200113
rect 194447 200085 194481 200113
rect 194509 200085 209779 200113
rect 209807 200085 209841 200113
rect 209869 200085 225139 200113
rect 225167 200085 225201 200113
rect 225229 200085 240499 200113
rect 240527 200085 240561 200113
rect 240589 200085 255859 200113
rect 255887 200085 255921 200113
rect 255949 200085 271219 200113
rect 271247 200085 271281 200113
rect 271309 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298990 200113
rect -958 200051 298990 200085
rect -958 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 33477 200051
rect 33505 200023 33539 200051
rect 33567 200023 33601 200051
rect 33629 200023 33663 200051
rect 33691 200023 48837 200051
rect 48865 200023 48899 200051
rect 48927 200023 48961 200051
rect 48989 200023 49023 200051
rect 49051 200023 64197 200051
rect 64225 200023 64259 200051
rect 64287 200023 64321 200051
rect 64349 200023 64383 200051
rect 64411 200023 79557 200051
rect 79585 200023 79619 200051
rect 79647 200023 79681 200051
rect 79709 200023 79743 200051
rect 79771 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 102259 200051
rect 102287 200023 102321 200051
rect 102349 200023 117619 200051
rect 117647 200023 117681 200051
rect 117709 200023 132979 200051
rect 133007 200023 133041 200051
rect 133069 200023 148339 200051
rect 148367 200023 148401 200051
rect 148429 200023 163699 200051
rect 163727 200023 163761 200051
rect 163789 200023 179059 200051
rect 179087 200023 179121 200051
rect 179149 200023 194419 200051
rect 194447 200023 194481 200051
rect 194509 200023 209779 200051
rect 209807 200023 209841 200051
rect 209869 200023 225139 200051
rect 225167 200023 225201 200051
rect 225229 200023 240499 200051
rect 240527 200023 240561 200051
rect 240589 200023 255859 200051
rect 255887 200023 255921 200051
rect 255949 200023 271219 200051
rect 271247 200023 271281 200051
rect 271309 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298990 200051
rect -958 199989 298990 200023
rect -958 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 33477 199989
rect 33505 199961 33539 199989
rect 33567 199961 33601 199989
rect 33629 199961 33663 199989
rect 33691 199961 48837 199989
rect 48865 199961 48899 199989
rect 48927 199961 48961 199989
rect 48989 199961 49023 199989
rect 49051 199961 64197 199989
rect 64225 199961 64259 199989
rect 64287 199961 64321 199989
rect 64349 199961 64383 199989
rect 64411 199961 79557 199989
rect 79585 199961 79619 199989
rect 79647 199961 79681 199989
rect 79709 199961 79743 199989
rect 79771 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 102259 199989
rect 102287 199961 102321 199989
rect 102349 199961 117619 199989
rect 117647 199961 117681 199989
rect 117709 199961 132979 199989
rect 133007 199961 133041 199989
rect 133069 199961 148339 199989
rect 148367 199961 148401 199989
rect 148429 199961 163699 199989
rect 163727 199961 163761 199989
rect 163789 199961 179059 199989
rect 179087 199961 179121 199989
rect 179149 199961 194419 199989
rect 194447 199961 194481 199989
rect 194509 199961 209779 199989
rect 209807 199961 209841 199989
rect 209869 199961 225139 199989
rect 225167 199961 225201 199989
rect 225229 199961 240499 199989
rect 240527 199961 240561 199989
rect 240589 199961 255859 199989
rect 255887 199961 255921 199989
rect 255949 199961 271219 199989
rect 271247 199961 271281 199989
rect 271309 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298990 199989
rect -958 199913 298990 199961
rect -958 194175 298990 194223
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 19977 194175
rect 20005 194147 20039 194175
rect 20067 194147 20101 194175
rect 20129 194147 20163 194175
rect 20191 194147 35337 194175
rect 35365 194147 35399 194175
rect 35427 194147 35461 194175
rect 35489 194147 35523 194175
rect 35551 194147 50697 194175
rect 50725 194147 50759 194175
rect 50787 194147 50821 194175
rect 50849 194147 50883 194175
rect 50911 194147 66057 194175
rect 66085 194147 66119 194175
rect 66147 194147 66181 194175
rect 66209 194147 66243 194175
rect 66271 194147 81417 194175
rect 81445 194147 81479 194175
rect 81507 194147 81541 194175
rect 81569 194147 81603 194175
rect 81631 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 109939 194175
rect 109967 194147 110001 194175
rect 110029 194147 125299 194175
rect 125327 194147 125361 194175
rect 125389 194147 140659 194175
rect 140687 194147 140721 194175
rect 140749 194147 156019 194175
rect 156047 194147 156081 194175
rect 156109 194147 171379 194175
rect 171407 194147 171441 194175
rect 171469 194147 186739 194175
rect 186767 194147 186801 194175
rect 186829 194147 202099 194175
rect 202127 194147 202161 194175
rect 202189 194147 217459 194175
rect 217487 194147 217521 194175
rect 217549 194147 232819 194175
rect 232847 194147 232881 194175
rect 232909 194147 248179 194175
rect 248207 194147 248241 194175
rect 248269 194147 263539 194175
rect 263567 194147 263601 194175
rect 263629 194147 278899 194175
rect 278927 194147 278961 194175
rect 278989 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect -958 194113 298990 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 19977 194113
rect 20005 194085 20039 194113
rect 20067 194085 20101 194113
rect 20129 194085 20163 194113
rect 20191 194085 35337 194113
rect 35365 194085 35399 194113
rect 35427 194085 35461 194113
rect 35489 194085 35523 194113
rect 35551 194085 50697 194113
rect 50725 194085 50759 194113
rect 50787 194085 50821 194113
rect 50849 194085 50883 194113
rect 50911 194085 66057 194113
rect 66085 194085 66119 194113
rect 66147 194085 66181 194113
rect 66209 194085 66243 194113
rect 66271 194085 81417 194113
rect 81445 194085 81479 194113
rect 81507 194085 81541 194113
rect 81569 194085 81603 194113
rect 81631 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 109939 194113
rect 109967 194085 110001 194113
rect 110029 194085 125299 194113
rect 125327 194085 125361 194113
rect 125389 194085 140659 194113
rect 140687 194085 140721 194113
rect 140749 194085 156019 194113
rect 156047 194085 156081 194113
rect 156109 194085 171379 194113
rect 171407 194085 171441 194113
rect 171469 194085 186739 194113
rect 186767 194085 186801 194113
rect 186829 194085 202099 194113
rect 202127 194085 202161 194113
rect 202189 194085 217459 194113
rect 217487 194085 217521 194113
rect 217549 194085 232819 194113
rect 232847 194085 232881 194113
rect 232909 194085 248179 194113
rect 248207 194085 248241 194113
rect 248269 194085 263539 194113
rect 263567 194085 263601 194113
rect 263629 194085 278899 194113
rect 278927 194085 278961 194113
rect 278989 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect -958 194051 298990 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 19977 194051
rect 20005 194023 20039 194051
rect 20067 194023 20101 194051
rect 20129 194023 20163 194051
rect 20191 194023 35337 194051
rect 35365 194023 35399 194051
rect 35427 194023 35461 194051
rect 35489 194023 35523 194051
rect 35551 194023 50697 194051
rect 50725 194023 50759 194051
rect 50787 194023 50821 194051
rect 50849 194023 50883 194051
rect 50911 194023 66057 194051
rect 66085 194023 66119 194051
rect 66147 194023 66181 194051
rect 66209 194023 66243 194051
rect 66271 194023 81417 194051
rect 81445 194023 81479 194051
rect 81507 194023 81541 194051
rect 81569 194023 81603 194051
rect 81631 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 109939 194051
rect 109967 194023 110001 194051
rect 110029 194023 125299 194051
rect 125327 194023 125361 194051
rect 125389 194023 140659 194051
rect 140687 194023 140721 194051
rect 140749 194023 156019 194051
rect 156047 194023 156081 194051
rect 156109 194023 171379 194051
rect 171407 194023 171441 194051
rect 171469 194023 186739 194051
rect 186767 194023 186801 194051
rect 186829 194023 202099 194051
rect 202127 194023 202161 194051
rect 202189 194023 217459 194051
rect 217487 194023 217521 194051
rect 217549 194023 232819 194051
rect 232847 194023 232881 194051
rect 232909 194023 248179 194051
rect 248207 194023 248241 194051
rect 248269 194023 263539 194051
rect 263567 194023 263601 194051
rect 263629 194023 278899 194051
rect 278927 194023 278961 194051
rect 278989 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect -958 193989 298990 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 19977 193989
rect 20005 193961 20039 193989
rect 20067 193961 20101 193989
rect 20129 193961 20163 193989
rect 20191 193961 35337 193989
rect 35365 193961 35399 193989
rect 35427 193961 35461 193989
rect 35489 193961 35523 193989
rect 35551 193961 50697 193989
rect 50725 193961 50759 193989
rect 50787 193961 50821 193989
rect 50849 193961 50883 193989
rect 50911 193961 66057 193989
rect 66085 193961 66119 193989
rect 66147 193961 66181 193989
rect 66209 193961 66243 193989
rect 66271 193961 81417 193989
rect 81445 193961 81479 193989
rect 81507 193961 81541 193989
rect 81569 193961 81603 193989
rect 81631 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 109939 193989
rect 109967 193961 110001 193989
rect 110029 193961 125299 193989
rect 125327 193961 125361 193989
rect 125389 193961 140659 193989
rect 140687 193961 140721 193989
rect 140749 193961 156019 193989
rect 156047 193961 156081 193989
rect 156109 193961 171379 193989
rect 171407 193961 171441 193989
rect 171469 193961 186739 193989
rect 186767 193961 186801 193989
rect 186829 193961 202099 193989
rect 202127 193961 202161 193989
rect 202189 193961 217459 193989
rect 217487 193961 217521 193989
rect 217549 193961 232819 193989
rect 232847 193961 232881 193989
rect 232909 193961 248179 193989
rect 248207 193961 248241 193989
rect 248269 193961 263539 193989
rect 263567 193961 263601 193989
rect 263629 193961 278899 193989
rect 278927 193961 278961 193989
rect 278989 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect -958 193913 298990 193961
rect -958 191175 298990 191223
rect -958 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 33477 191175
rect 33505 191147 33539 191175
rect 33567 191147 33601 191175
rect 33629 191147 33663 191175
rect 33691 191147 48837 191175
rect 48865 191147 48899 191175
rect 48927 191147 48961 191175
rect 48989 191147 49023 191175
rect 49051 191147 64197 191175
rect 64225 191147 64259 191175
rect 64287 191147 64321 191175
rect 64349 191147 64383 191175
rect 64411 191147 79557 191175
rect 79585 191147 79619 191175
rect 79647 191147 79681 191175
rect 79709 191147 79743 191175
rect 79771 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 102259 191175
rect 102287 191147 102321 191175
rect 102349 191147 117619 191175
rect 117647 191147 117681 191175
rect 117709 191147 132979 191175
rect 133007 191147 133041 191175
rect 133069 191147 148339 191175
rect 148367 191147 148401 191175
rect 148429 191147 163699 191175
rect 163727 191147 163761 191175
rect 163789 191147 179059 191175
rect 179087 191147 179121 191175
rect 179149 191147 194419 191175
rect 194447 191147 194481 191175
rect 194509 191147 209779 191175
rect 209807 191147 209841 191175
rect 209869 191147 225139 191175
rect 225167 191147 225201 191175
rect 225229 191147 240499 191175
rect 240527 191147 240561 191175
rect 240589 191147 255859 191175
rect 255887 191147 255921 191175
rect 255949 191147 271219 191175
rect 271247 191147 271281 191175
rect 271309 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298990 191175
rect -958 191113 298990 191147
rect -958 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 33477 191113
rect 33505 191085 33539 191113
rect 33567 191085 33601 191113
rect 33629 191085 33663 191113
rect 33691 191085 48837 191113
rect 48865 191085 48899 191113
rect 48927 191085 48961 191113
rect 48989 191085 49023 191113
rect 49051 191085 64197 191113
rect 64225 191085 64259 191113
rect 64287 191085 64321 191113
rect 64349 191085 64383 191113
rect 64411 191085 79557 191113
rect 79585 191085 79619 191113
rect 79647 191085 79681 191113
rect 79709 191085 79743 191113
rect 79771 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 102259 191113
rect 102287 191085 102321 191113
rect 102349 191085 117619 191113
rect 117647 191085 117681 191113
rect 117709 191085 132979 191113
rect 133007 191085 133041 191113
rect 133069 191085 148339 191113
rect 148367 191085 148401 191113
rect 148429 191085 163699 191113
rect 163727 191085 163761 191113
rect 163789 191085 179059 191113
rect 179087 191085 179121 191113
rect 179149 191085 194419 191113
rect 194447 191085 194481 191113
rect 194509 191085 209779 191113
rect 209807 191085 209841 191113
rect 209869 191085 225139 191113
rect 225167 191085 225201 191113
rect 225229 191085 240499 191113
rect 240527 191085 240561 191113
rect 240589 191085 255859 191113
rect 255887 191085 255921 191113
rect 255949 191085 271219 191113
rect 271247 191085 271281 191113
rect 271309 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298990 191113
rect -958 191051 298990 191085
rect -958 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 33477 191051
rect 33505 191023 33539 191051
rect 33567 191023 33601 191051
rect 33629 191023 33663 191051
rect 33691 191023 48837 191051
rect 48865 191023 48899 191051
rect 48927 191023 48961 191051
rect 48989 191023 49023 191051
rect 49051 191023 64197 191051
rect 64225 191023 64259 191051
rect 64287 191023 64321 191051
rect 64349 191023 64383 191051
rect 64411 191023 79557 191051
rect 79585 191023 79619 191051
rect 79647 191023 79681 191051
rect 79709 191023 79743 191051
rect 79771 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 102259 191051
rect 102287 191023 102321 191051
rect 102349 191023 117619 191051
rect 117647 191023 117681 191051
rect 117709 191023 132979 191051
rect 133007 191023 133041 191051
rect 133069 191023 148339 191051
rect 148367 191023 148401 191051
rect 148429 191023 163699 191051
rect 163727 191023 163761 191051
rect 163789 191023 179059 191051
rect 179087 191023 179121 191051
rect 179149 191023 194419 191051
rect 194447 191023 194481 191051
rect 194509 191023 209779 191051
rect 209807 191023 209841 191051
rect 209869 191023 225139 191051
rect 225167 191023 225201 191051
rect 225229 191023 240499 191051
rect 240527 191023 240561 191051
rect 240589 191023 255859 191051
rect 255887 191023 255921 191051
rect 255949 191023 271219 191051
rect 271247 191023 271281 191051
rect 271309 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298990 191051
rect -958 190989 298990 191023
rect -958 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 33477 190989
rect 33505 190961 33539 190989
rect 33567 190961 33601 190989
rect 33629 190961 33663 190989
rect 33691 190961 48837 190989
rect 48865 190961 48899 190989
rect 48927 190961 48961 190989
rect 48989 190961 49023 190989
rect 49051 190961 64197 190989
rect 64225 190961 64259 190989
rect 64287 190961 64321 190989
rect 64349 190961 64383 190989
rect 64411 190961 79557 190989
rect 79585 190961 79619 190989
rect 79647 190961 79681 190989
rect 79709 190961 79743 190989
rect 79771 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 102259 190989
rect 102287 190961 102321 190989
rect 102349 190961 117619 190989
rect 117647 190961 117681 190989
rect 117709 190961 132979 190989
rect 133007 190961 133041 190989
rect 133069 190961 148339 190989
rect 148367 190961 148401 190989
rect 148429 190961 163699 190989
rect 163727 190961 163761 190989
rect 163789 190961 179059 190989
rect 179087 190961 179121 190989
rect 179149 190961 194419 190989
rect 194447 190961 194481 190989
rect 194509 190961 209779 190989
rect 209807 190961 209841 190989
rect 209869 190961 225139 190989
rect 225167 190961 225201 190989
rect 225229 190961 240499 190989
rect 240527 190961 240561 190989
rect 240589 190961 255859 190989
rect 255887 190961 255921 190989
rect 255949 190961 271219 190989
rect 271247 190961 271281 190989
rect 271309 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298990 190989
rect -958 190913 298990 190961
rect -958 185175 298990 185223
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 19977 185175
rect 20005 185147 20039 185175
rect 20067 185147 20101 185175
rect 20129 185147 20163 185175
rect 20191 185147 35337 185175
rect 35365 185147 35399 185175
rect 35427 185147 35461 185175
rect 35489 185147 35523 185175
rect 35551 185147 50697 185175
rect 50725 185147 50759 185175
rect 50787 185147 50821 185175
rect 50849 185147 50883 185175
rect 50911 185147 66057 185175
rect 66085 185147 66119 185175
rect 66147 185147 66181 185175
rect 66209 185147 66243 185175
rect 66271 185147 81417 185175
rect 81445 185147 81479 185175
rect 81507 185147 81541 185175
rect 81569 185147 81603 185175
rect 81631 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 109939 185175
rect 109967 185147 110001 185175
rect 110029 185147 125299 185175
rect 125327 185147 125361 185175
rect 125389 185147 140659 185175
rect 140687 185147 140721 185175
rect 140749 185147 156019 185175
rect 156047 185147 156081 185175
rect 156109 185147 171379 185175
rect 171407 185147 171441 185175
rect 171469 185147 186739 185175
rect 186767 185147 186801 185175
rect 186829 185147 202099 185175
rect 202127 185147 202161 185175
rect 202189 185147 217459 185175
rect 217487 185147 217521 185175
rect 217549 185147 232819 185175
rect 232847 185147 232881 185175
rect 232909 185147 248179 185175
rect 248207 185147 248241 185175
rect 248269 185147 263539 185175
rect 263567 185147 263601 185175
rect 263629 185147 278899 185175
rect 278927 185147 278961 185175
rect 278989 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect -958 185113 298990 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 19977 185113
rect 20005 185085 20039 185113
rect 20067 185085 20101 185113
rect 20129 185085 20163 185113
rect 20191 185085 35337 185113
rect 35365 185085 35399 185113
rect 35427 185085 35461 185113
rect 35489 185085 35523 185113
rect 35551 185085 50697 185113
rect 50725 185085 50759 185113
rect 50787 185085 50821 185113
rect 50849 185085 50883 185113
rect 50911 185085 66057 185113
rect 66085 185085 66119 185113
rect 66147 185085 66181 185113
rect 66209 185085 66243 185113
rect 66271 185085 81417 185113
rect 81445 185085 81479 185113
rect 81507 185085 81541 185113
rect 81569 185085 81603 185113
rect 81631 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 109939 185113
rect 109967 185085 110001 185113
rect 110029 185085 125299 185113
rect 125327 185085 125361 185113
rect 125389 185085 140659 185113
rect 140687 185085 140721 185113
rect 140749 185085 156019 185113
rect 156047 185085 156081 185113
rect 156109 185085 171379 185113
rect 171407 185085 171441 185113
rect 171469 185085 186739 185113
rect 186767 185085 186801 185113
rect 186829 185085 202099 185113
rect 202127 185085 202161 185113
rect 202189 185085 217459 185113
rect 217487 185085 217521 185113
rect 217549 185085 232819 185113
rect 232847 185085 232881 185113
rect 232909 185085 248179 185113
rect 248207 185085 248241 185113
rect 248269 185085 263539 185113
rect 263567 185085 263601 185113
rect 263629 185085 278899 185113
rect 278927 185085 278961 185113
rect 278989 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect -958 185051 298990 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 19977 185051
rect 20005 185023 20039 185051
rect 20067 185023 20101 185051
rect 20129 185023 20163 185051
rect 20191 185023 35337 185051
rect 35365 185023 35399 185051
rect 35427 185023 35461 185051
rect 35489 185023 35523 185051
rect 35551 185023 50697 185051
rect 50725 185023 50759 185051
rect 50787 185023 50821 185051
rect 50849 185023 50883 185051
rect 50911 185023 66057 185051
rect 66085 185023 66119 185051
rect 66147 185023 66181 185051
rect 66209 185023 66243 185051
rect 66271 185023 81417 185051
rect 81445 185023 81479 185051
rect 81507 185023 81541 185051
rect 81569 185023 81603 185051
rect 81631 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 109939 185051
rect 109967 185023 110001 185051
rect 110029 185023 125299 185051
rect 125327 185023 125361 185051
rect 125389 185023 140659 185051
rect 140687 185023 140721 185051
rect 140749 185023 156019 185051
rect 156047 185023 156081 185051
rect 156109 185023 171379 185051
rect 171407 185023 171441 185051
rect 171469 185023 186739 185051
rect 186767 185023 186801 185051
rect 186829 185023 202099 185051
rect 202127 185023 202161 185051
rect 202189 185023 217459 185051
rect 217487 185023 217521 185051
rect 217549 185023 232819 185051
rect 232847 185023 232881 185051
rect 232909 185023 248179 185051
rect 248207 185023 248241 185051
rect 248269 185023 263539 185051
rect 263567 185023 263601 185051
rect 263629 185023 278899 185051
rect 278927 185023 278961 185051
rect 278989 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect -958 184989 298990 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 19977 184989
rect 20005 184961 20039 184989
rect 20067 184961 20101 184989
rect 20129 184961 20163 184989
rect 20191 184961 35337 184989
rect 35365 184961 35399 184989
rect 35427 184961 35461 184989
rect 35489 184961 35523 184989
rect 35551 184961 50697 184989
rect 50725 184961 50759 184989
rect 50787 184961 50821 184989
rect 50849 184961 50883 184989
rect 50911 184961 66057 184989
rect 66085 184961 66119 184989
rect 66147 184961 66181 184989
rect 66209 184961 66243 184989
rect 66271 184961 81417 184989
rect 81445 184961 81479 184989
rect 81507 184961 81541 184989
rect 81569 184961 81603 184989
rect 81631 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 109939 184989
rect 109967 184961 110001 184989
rect 110029 184961 125299 184989
rect 125327 184961 125361 184989
rect 125389 184961 140659 184989
rect 140687 184961 140721 184989
rect 140749 184961 156019 184989
rect 156047 184961 156081 184989
rect 156109 184961 171379 184989
rect 171407 184961 171441 184989
rect 171469 184961 186739 184989
rect 186767 184961 186801 184989
rect 186829 184961 202099 184989
rect 202127 184961 202161 184989
rect 202189 184961 217459 184989
rect 217487 184961 217521 184989
rect 217549 184961 232819 184989
rect 232847 184961 232881 184989
rect 232909 184961 248179 184989
rect 248207 184961 248241 184989
rect 248269 184961 263539 184989
rect 263567 184961 263601 184989
rect 263629 184961 278899 184989
rect 278927 184961 278961 184989
rect 278989 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect -958 184913 298990 184961
rect -958 182175 298990 182223
rect -958 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 33477 182175
rect 33505 182147 33539 182175
rect 33567 182147 33601 182175
rect 33629 182147 33663 182175
rect 33691 182147 48837 182175
rect 48865 182147 48899 182175
rect 48927 182147 48961 182175
rect 48989 182147 49023 182175
rect 49051 182147 64197 182175
rect 64225 182147 64259 182175
rect 64287 182147 64321 182175
rect 64349 182147 64383 182175
rect 64411 182147 79557 182175
rect 79585 182147 79619 182175
rect 79647 182147 79681 182175
rect 79709 182147 79743 182175
rect 79771 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 102259 182175
rect 102287 182147 102321 182175
rect 102349 182147 117619 182175
rect 117647 182147 117681 182175
rect 117709 182147 132979 182175
rect 133007 182147 133041 182175
rect 133069 182147 148339 182175
rect 148367 182147 148401 182175
rect 148429 182147 163699 182175
rect 163727 182147 163761 182175
rect 163789 182147 179059 182175
rect 179087 182147 179121 182175
rect 179149 182147 194419 182175
rect 194447 182147 194481 182175
rect 194509 182147 209779 182175
rect 209807 182147 209841 182175
rect 209869 182147 225139 182175
rect 225167 182147 225201 182175
rect 225229 182147 240499 182175
rect 240527 182147 240561 182175
rect 240589 182147 255859 182175
rect 255887 182147 255921 182175
rect 255949 182147 271219 182175
rect 271247 182147 271281 182175
rect 271309 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298990 182175
rect -958 182113 298990 182147
rect -958 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 33477 182113
rect 33505 182085 33539 182113
rect 33567 182085 33601 182113
rect 33629 182085 33663 182113
rect 33691 182085 48837 182113
rect 48865 182085 48899 182113
rect 48927 182085 48961 182113
rect 48989 182085 49023 182113
rect 49051 182085 64197 182113
rect 64225 182085 64259 182113
rect 64287 182085 64321 182113
rect 64349 182085 64383 182113
rect 64411 182085 79557 182113
rect 79585 182085 79619 182113
rect 79647 182085 79681 182113
rect 79709 182085 79743 182113
rect 79771 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 102259 182113
rect 102287 182085 102321 182113
rect 102349 182085 117619 182113
rect 117647 182085 117681 182113
rect 117709 182085 132979 182113
rect 133007 182085 133041 182113
rect 133069 182085 148339 182113
rect 148367 182085 148401 182113
rect 148429 182085 163699 182113
rect 163727 182085 163761 182113
rect 163789 182085 179059 182113
rect 179087 182085 179121 182113
rect 179149 182085 194419 182113
rect 194447 182085 194481 182113
rect 194509 182085 209779 182113
rect 209807 182085 209841 182113
rect 209869 182085 225139 182113
rect 225167 182085 225201 182113
rect 225229 182085 240499 182113
rect 240527 182085 240561 182113
rect 240589 182085 255859 182113
rect 255887 182085 255921 182113
rect 255949 182085 271219 182113
rect 271247 182085 271281 182113
rect 271309 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298990 182113
rect -958 182051 298990 182085
rect -958 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 33477 182051
rect 33505 182023 33539 182051
rect 33567 182023 33601 182051
rect 33629 182023 33663 182051
rect 33691 182023 48837 182051
rect 48865 182023 48899 182051
rect 48927 182023 48961 182051
rect 48989 182023 49023 182051
rect 49051 182023 64197 182051
rect 64225 182023 64259 182051
rect 64287 182023 64321 182051
rect 64349 182023 64383 182051
rect 64411 182023 79557 182051
rect 79585 182023 79619 182051
rect 79647 182023 79681 182051
rect 79709 182023 79743 182051
rect 79771 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 102259 182051
rect 102287 182023 102321 182051
rect 102349 182023 117619 182051
rect 117647 182023 117681 182051
rect 117709 182023 132979 182051
rect 133007 182023 133041 182051
rect 133069 182023 148339 182051
rect 148367 182023 148401 182051
rect 148429 182023 163699 182051
rect 163727 182023 163761 182051
rect 163789 182023 179059 182051
rect 179087 182023 179121 182051
rect 179149 182023 194419 182051
rect 194447 182023 194481 182051
rect 194509 182023 209779 182051
rect 209807 182023 209841 182051
rect 209869 182023 225139 182051
rect 225167 182023 225201 182051
rect 225229 182023 240499 182051
rect 240527 182023 240561 182051
rect 240589 182023 255859 182051
rect 255887 182023 255921 182051
rect 255949 182023 271219 182051
rect 271247 182023 271281 182051
rect 271309 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298990 182051
rect -958 181989 298990 182023
rect -958 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 33477 181989
rect 33505 181961 33539 181989
rect 33567 181961 33601 181989
rect 33629 181961 33663 181989
rect 33691 181961 48837 181989
rect 48865 181961 48899 181989
rect 48927 181961 48961 181989
rect 48989 181961 49023 181989
rect 49051 181961 64197 181989
rect 64225 181961 64259 181989
rect 64287 181961 64321 181989
rect 64349 181961 64383 181989
rect 64411 181961 79557 181989
rect 79585 181961 79619 181989
rect 79647 181961 79681 181989
rect 79709 181961 79743 181989
rect 79771 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 102259 181989
rect 102287 181961 102321 181989
rect 102349 181961 117619 181989
rect 117647 181961 117681 181989
rect 117709 181961 132979 181989
rect 133007 181961 133041 181989
rect 133069 181961 148339 181989
rect 148367 181961 148401 181989
rect 148429 181961 163699 181989
rect 163727 181961 163761 181989
rect 163789 181961 179059 181989
rect 179087 181961 179121 181989
rect 179149 181961 194419 181989
rect 194447 181961 194481 181989
rect 194509 181961 209779 181989
rect 209807 181961 209841 181989
rect 209869 181961 225139 181989
rect 225167 181961 225201 181989
rect 225229 181961 240499 181989
rect 240527 181961 240561 181989
rect 240589 181961 255859 181989
rect 255887 181961 255921 181989
rect 255949 181961 271219 181989
rect 271247 181961 271281 181989
rect 271309 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298990 181989
rect -958 181913 298990 181961
rect -958 176175 298990 176223
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 19977 176175
rect 20005 176147 20039 176175
rect 20067 176147 20101 176175
rect 20129 176147 20163 176175
rect 20191 176147 35337 176175
rect 35365 176147 35399 176175
rect 35427 176147 35461 176175
rect 35489 176147 35523 176175
rect 35551 176147 50697 176175
rect 50725 176147 50759 176175
rect 50787 176147 50821 176175
rect 50849 176147 50883 176175
rect 50911 176147 66057 176175
rect 66085 176147 66119 176175
rect 66147 176147 66181 176175
rect 66209 176147 66243 176175
rect 66271 176147 81417 176175
rect 81445 176147 81479 176175
rect 81507 176147 81541 176175
rect 81569 176147 81603 176175
rect 81631 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 109939 176175
rect 109967 176147 110001 176175
rect 110029 176147 125299 176175
rect 125327 176147 125361 176175
rect 125389 176147 140659 176175
rect 140687 176147 140721 176175
rect 140749 176147 156019 176175
rect 156047 176147 156081 176175
rect 156109 176147 171379 176175
rect 171407 176147 171441 176175
rect 171469 176147 186739 176175
rect 186767 176147 186801 176175
rect 186829 176147 202099 176175
rect 202127 176147 202161 176175
rect 202189 176147 217459 176175
rect 217487 176147 217521 176175
rect 217549 176147 232819 176175
rect 232847 176147 232881 176175
rect 232909 176147 248179 176175
rect 248207 176147 248241 176175
rect 248269 176147 263539 176175
rect 263567 176147 263601 176175
rect 263629 176147 278899 176175
rect 278927 176147 278961 176175
rect 278989 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect -958 176113 298990 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 19977 176113
rect 20005 176085 20039 176113
rect 20067 176085 20101 176113
rect 20129 176085 20163 176113
rect 20191 176085 35337 176113
rect 35365 176085 35399 176113
rect 35427 176085 35461 176113
rect 35489 176085 35523 176113
rect 35551 176085 50697 176113
rect 50725 176085 50759 176113
rect 50787 176085 50821 176113
rect 50849 176085 50883 176113
rect 50911 176085 66057 176113
rect 66085 176085 66119 176113
rect 66147 176085 66181 176113
rect 66209 176085 66243 176113
rect 66271 176085 81417 176113
rect 81445 176085 81479 176113
rect 81507 176085 81541 176113
rect 81569 176085 81603 176113
rect 81631 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 109939 176113
rect 109967 176085 110001 176113
rect 110029 176085 125299 176113
rect 125327 176085 125361 176113
rect 125389 176085 140659 176113
rect 140687 176085 140721 176113
rect 140749 176085 156019 176113
rect 156047 176085 156081 176113
rect 156109 176085 171379 176113
rect 171407 176085 171441 176113
rect 171469 176085 186739 176113
rect 186767 176085 186801 176113
rect 186829 176085 202099 176113
rect 202127 176085 202161 176113
rect 202189 176085 217459 176113
rect 217487 176085 217521 176113
rect 217549 176085 232819 176113
rect 232847 176085 232881 176113
rect 232909 176085 248179 176113
rect 248207 176085 248241 176113
rect 248269 176085 263539 176113
rect 263567 176085 263601 176113
rect 263629 176085 278899 176113
rect 278927 176085 278961 176113
rect 278989 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect -958 176051 298990 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 19977 176051
rect 20005 176023 20039 176051
rect 20067 176023 20101 176051
rect 20129 176023 20163 176051
rect 20191 176023 35337 176051
rect 35365 176023 35399 176051
rect 35427 176023 35461 176051
rect 35489 176023 35523 176051
rect 35551 176023 50697 176051
rect 50725 176023 50759 176051
rect 50787 176023 50821 176051
rect 50849 176023 50883 176051
rect 50911 176023 66057 176051
rect 66085 176023 66119 176051
rect 66147 176023 66181 176051
rect 66209 176023 66243 176051
rect 66271 176023 81417 176051
rect 81445 176023 81479 176051
rect 81507 176023 81541 176051
rect 81569 176023 81603 176051
rect 81631 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 109939 176051
rect 109967 176023 110001 176051
rect 110029 176023 125299 176051
rect 125327 176023 125361 176051
rect 125389 176023 140659 176051
rect 140687 176023 140721 176051
rect 140749 176023 156019 176051
rect 156047 176023 156081 176051
rect 156109 176023 171379 176051
rect 171407 176023 171441 176051
rect 171469 176023 186739 176051
rect 186767 176023 186801 176051
rect 186829 176023 202099 176051
rect 202127 176023 202161 176051
rect 202189 176023 217459 176051
rect 217487 176023 217521 176051
rect 217549 176023 232819 176051
rect 232847 176023 232881 176051
rect 232909 176023 248179 176051
rect 248207 176023 248241 176051
rect 248269 176023 263539 176051
rect 263567 176023 263601 176051
rect 263629 176023 278899 176051
rect 278927 176023 278961 176051
rect 278989 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect -958 175989 298990 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 19977 175989
rect 20005 175961 20039 175989
rect 20067 175961 20101 175989
rect 20129 175961 20163 175989
rect 20191 175961 35337 175989
rect 35365 175961 35399 175989
rect 35427 175961 35461 175989
rect 35489 175961 35523 175989
rect 35551 175961 50697 175989
rect 50725 175961 50759 175989
rect 50787 175961 50821 175989
rect 50849 175961 50883 175989
rect 50911 175961 66057 175989
rect 66085 175961 66119 175989
rect 66147 175961 66181 175989
rect 66209 175961 66243 175989
rect 66271 175961 81417 175989
rect 81445 175961 81479 175989
rect 81507 175961 81541 175989
rect 81569 175961 81603 175989
rect 81631 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 109939 175989
rect 109967 175961 110001 175989
rect 110029 175961 125299 175989
rect 125327 175961 125361 175989
rect 125389 175961 140659 175989
rect 140687 175961 140721 175989
rect 140749 175961 156019 175989
rect 156047 175961 156081 175989
rect 156109 175961 171379 175989
rect 171407 175961 171441 175989
rect 171469 175961 186739 175989
rect 186767 175961 186801 175989
rect 186829 175961 202099 175989
rect 202127 175961 202161 175989
rect 202189 175961 217459 175989
rect 217487 175961 217521 175989
rect 217549 175961 232819 175989
rect 232847 175961 232881 175989
rect 232909 175961 248179 175989
rect 248207 175961 248241 175989
rect 248269 175961 263539 175989
rect 263567 175961 263601 175989
rect 263629 175961 278899 175989
rect 278927 175961 278961 175989
rect 278989 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect -958 175913 298990 175961
rect -958 173175 298990 173223
rect -958 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 33477 173175
rect 33505 173147 33539 173175
rect 33567 173147 33601 173175
rect 33629 173147 33663 173175
rect 33691 173147 48837 173175
rect 48865 173147 48899 173175
rect 48927 173147 48961 173175
rect 48989 173147 49023 173175
rect 49051 173147 64197 173175
rect 64225 173147 64259 173175
rect 64287 173147 64321 173175
rect 64349 173147 64383 173175
rect 64411 173147 79557 173175
rect 79585 173147 79619 173175
rect 79647 173147 79681 173175
rect 79709 173147 79743 173175
rect 79771 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 102259 173175
rect 102287 173147 102321 173175
rect 102349 173147 117619 173175
rect 117647 173147 117681 173175
rect 117709 173147 132979 173175
rect 133007 173147 133041 173175
rect 133069 173147 148339 173175
rect 148367 173147 148401 173175
rect 148429 173147 163699 173175
rect 163727 173147 163761 173175
rect 163789 173147 179059 173175
rect 179087 173147 179121 173175
rect 179149 173147 194419 173175
rect 194447 173147 194481 173175
rect 194509 173147 209779 173175
rect 209807 173147 209841 173175
rect 209869 173147 225139 173175
rect 225167 173147 225201 173175
rect 225229 173147 240499 173175
rect 240527 173147 240561 173175
rect 240589 173147 255859 173175
rect 255887 173147 255921 173175
rect 255949 173147 271219 173175
rect 271247 173147 271281 173175
rect 271309 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298990 173175
rect -958 173113 298990 173147
rect -958 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 33477 173113
rect 33505 173085 33539 173113
rect 33567 173085 33601 173113
rect 33629 173085 33663 173113
rect 33691 173085 48837 173113
rect 48865 173085 48899 173113
rect 48927 173085 48961 173113
rect 48989 173085 49023 173113
rect 49051 173085 64197 173113
rect 64225 173085 64259 173113
rect 64287 173085 64321 173113
rect 64349 173085 64383 173113
rect 64411 173085 79557 173113
rect 79585 173085 79619 173113
rect 79647 173085 79681 173113
rect 79709 173085 79743 173113
rect 79771 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 102259 173113
rect 102287 173085 102321 173113
rect 102349 173085 117619 173113
rect 117647 173085 117681 173113
rect 117709 173085 132979 173113
rect 133007 173085 133041 173113
rect 133069 173085 148339 173113
rect 148367 173085 148401 173113
rect 148429 173085 163699 173113
rect 163727 173085 163761 173113
rect 163789 173085 179059 173113
rect 179087 173085 179121 173113
rect 179149 173085 194419 173113
rect 194447 173085 194481 173113
rect 194509 173085 209779 173113
rect 209807 173085 209841 173113
rect 209869 173085 225139 173113
rect 225167 173085 225201 173113
rect 225229 173085 240499 173113
rect 240527 173085 240561 173113
rect 240589 173085 255859 173113
rect 255887 173085 255921 173113
rect 255949 173085 271219 173113
rect 271247 173085 271281 173113
rect 271309 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298990 173113
rect -958 173051 298990 173085
rect -958 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 33477 173051
rect 33505 173023 33539 173051
rect 33567 173023 33601 173051
rect 33629 173023 33663 173051
rect 33691 173023 48837 173051
rect 48865 173023 48899 173051
rect 48927 173023 48961 173051
rect 48989 173023 49023 173051
rect 49051 173023 64197 173051
rect 64225 173023 64259 173051
rect 64287 173023 64321 173051
rect 64349 173023 64383 173051
rect 64411 173023 79557 173051
rect 79585 173023 79619 173051
rect 79647 173023 79681 173051
rect 79709 173023 79743 173051
rect 79771 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 102259 173051
rect 102287 173023 102321 173051
rect 102349 173023 117619 173051
rect 117647 173023 117681 173051
rect 117709 173023 132979 173051
rect 133007 173023 133041 173051
rect 133069 173023 148339 173051
rect 148367 173023 148401 173051
rect 148429 173023 163699 173051
rect 163727 173023 163761 173051
rect 163789 173023 179059 173051
rect 179087 173023 179121 173051
rect 179149 173023 194419 173051
rect 194447 173023 194481 173051
rect 194509 173023 209779 173051
rect 209807 173023 209841 173051
rect 209869 173023 225139 173051
rect 225167 173023 225201 173051
rect 225229 173023 240499 173051
rect 240527 173023 240561 173051
rect 240589 173023 255859 173051
rect 255887 173023 255921 173051
rect 255949 173023 271219 173051
rect 271247 173023 271281 173051
rect 271309 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298990 173051
rect -958 172989 298990 173023
rect -958 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 33477 172989
rect 33505 172961 33539 172989
rect 33567 172961 33601 172989
rect 33629 172961 33663 172989
rect 33691 172961 48837 172989
rect 48865 172961 48899 172989
rect 48927 172961 48961 172989
rect 48989 172961 49023 172989
rect 49051 172961 64197 172989
rect 64225 172961 64259 172989
rect 64287 172961 64321 172989
rect 64349 172961 64383 172989
rect 64411 172961 79557 172989
rect 79585 172961 79619 172989
rect 79647 172961 79681 172989
rect 79709 172961 79743 172989
rect 79771 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 102259 172989
rect 102287 172961 102321 172989
rect 102349 172961 117619 172989
rect 117647 172961 117681 172989
rect 117709 172961 132979 172989
rect 133007 172961 133041 172989
rect 133069 172961 148339 172989
rect 148367 172961 148401 172989
rect 148429 172961 163699 172989
rect 163727 172961 163761 172989
rect 163789 172961 179059 172989
rect 179087 172961 179121 172989
rect 179149 172961 194419 172989
rect 194447 172961 194481 172989
rect 194509 172961 209779 172989
rect 209807 172961 209841 172989
rect 209869 172961 225139 172989
rect 225167 172961 225201 172989
rect 225229 172961 240499 172989
rect 240527 172961 240561 172989
rect 240589 172961 255859 172989
rect 255887 172961 255921 172989
rect 255949 172961 271219 172989
rect 271247 172961 271281 172989
rect 271309 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298990 172989
rect -958 172913 298990 172961
rect -958 167175 298990 167223
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 109939 167175
rect 109967 167147 110001 167175
rect 110029 167147 125299 167175
rect 125327 167147 125361 167175
rect 125389 167147 140659 167175
rect 140687 167147 140721 167175
rect 140749 167147 156019 167175
rect 156047 167147 156081 167175
rect 156109 167147 171379 167175
rect 171407 167147 171441 167175
rect 171469 167147 186739 167175
rect 186767 167147 186801 167175
rect 186829 167147 202099 167175
rect 202127 167147 202161 167175
rect 202189 167147 217459 167175
rect 217487 167147 217521 167175
rect 217549 167147 232819 167175
rect 232847 167147 232881 167175
rect 232909 167147 248179 167175
rect 248207 167147 248241 167175
rect 248269 167147 263539 167175
rect 263567 167147 263601 167175
rect 263629 167147 278899 167175
rect 278927 167147 278961 167175
rect 278989 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect -958 167113 298990 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 109939 167113
rect 109967 167085 110001 167113
rect 110029 167085 125299 167113
rect 125327 167085 125361 167113
rect 125389 167085 140659 167113
rect 140687 167085 140721 167113
rect 140749 167085 156019 167113
rect 156047 167085 156081 167113
rect 156109 167085 171379 167113
rect 171407 167085 171441 167113
rect 171469 167085 186739 167113
rect 186767 167085 186801 167113
rect 186829 167085 202099 167113
rect 202127 167085 202161 167113
rect 202189 167085 217459 167113
rect 217487 167085 217521 167113
rect 217549 167085 232819 167113
rect 232847 167085 232881 167113
rect 232909 167085 248179 167113
rect 248207 167085 248241 167113
rect 248269 167085 263539 167113
rect 263567 167085 263601 167113
rect 263629 167085 278899 167113
rect 278927 167085 278961 167113
rect 278989 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect -958 167051 298990 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 109939 167051
rect 109967 167023 110001 167051
rect 110029 167023 125299 167051
rect 125327 167023 125361 167051
rect 125389 167023 140659 167051
rect 140687 167023 140721 167051
rect 140749 167023 156019 167051
rect 156047 167023 156081 167051
rect 156109 167023 171379 167051
rect 171407 167023 171441 167051
rect 171469 167023 186739 167051
rect 186767 167023 186801 167051
rect 186829 167023 202099 167051
rect 202127 167023 202161 167051
rect 202189 167023 217459 167051
rect 217487 167023 217521 167051
rect 217549 167023 232819 167051
rect 232847 167023 232881 167051
rect 232909 167023 248179 167051
rect 248207 167023 248241 167051
rect 248269 167023 263539 167051
rect 263567 167023 263601 167051
rect 263629 167023 278899 167051
rect 278927 167023 278961 167051
rect 278989 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect -958 166989 298990 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 109939 166989
rect 109967 166961 110001 166989
rect 110029 166961 125299 166989
rect 125327 166961 125361 166989
rect 125389 166961 140659 166989
rect 140687 166961 140721 166989
rect 140749 166961 156019 166989
rect 156047 166961 156081 166989
rect 156109 166961 171379 166989
rect 171407 166961 171441 166989
rect 171469 166961 186739 166989
rect 186767 166961 186801 166989
rect 186829 166961 202099 166989
rect 202127 166961 202161 166989
rect 202189 166961 217459 166989
rect 217487 166961 217521 166989
rect 217549 166961 232819 166989
rect 232847 166961 232881 166989
rect 232909 166961 248179 166989
rect 248207 166961 248241 166989
rect 248269 166961 263539 166989
rect 263567 166961 263601 166989
rect 263629 166961 278899 166989
rect 278927 166961 278961 166989
rect 278989 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect -958 166913 298990 166961
rect -958 164175 298990 164223
rect -958 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 102259 164175
rect 102287 164147 102321 164175
rect 102349 164147 117619 164175
rect 117647 164147 117681 164175
rect 117709 164147 132979 164175
rect 133007 164147 133041 164175
rect 133069 164147 148339 164175
rect 148367 164147 148401 164175
rect 148429 164147 163699 164175
rect 163727 164147 163761 164175
rect 163789 164147 179059 164175
rect 179087 164147 179121 164175
rect 179149 164147 194419 164175
rect 194447 164147 194481 164175
rect 194509 164147 209779 164175
rect 209807 164147 209841 164175
rect 209869 164147 225139 164175
rect 225167 164147 225201 164175
rect 225229 164147 240499 164175
rect 240527 164147 240561 164175
rect 240589 164147 255859 164175
rect 255887 164147 255921 164175
rect 255949 164147 271219 164175
rect 271247 164147 271281 164175
rect 271309 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298990 164175
rect -958 164113 298990 164147
rect -958 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 102259 164113
rect 102287 164085 102321 164113
rect 102349 164085 117619 164113
rect 117647 164085 117681 164113
rect 117709 164085 132979 164113
rect 133007 164085 133041 164113
rect 133069 164085 148339 164113
rect 148367 164085 148401 164113
rect 148429 164085 163699 164113
rect 163727 164085 163761 164113
rect 163789 164085 179059 164113
rect 179087 164085 179121 164113
rect 179149 164085 194419 164113
rect 194447 164085 194481 164113
rect 194509 164085 209779 164113
rect 209807 164085 209841 164113
rect 209869 164085 225139 164113
rect 225167 164085 225201 164113
rect 225229 164085 240499 164113
rect 240527 164085 240561 164113
rect 240589 164085 255859 164113
rect 255887 164085 255921 164113
rect 255949 164085 271219 164113
rect 271247 164085 271281 164113
rect 271309 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298990 164113
rect -958 164051 298990 164085
rect -958 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 102259 164051
rect 102287 164023 102321 164051
rect 102349 164023 117619 164051
rect 117647 164023 117681 164051
rect 117709 164023 132979 164051
rect 133007 164023 133041 164051
rect 133069 164023 148339 164051
rect 148367 164023 148401 164051
rect 148429 164023 163699 164051
rect 163727 164023 163761 164051
rect 163789 164023 179059 164051
rect 179087 164023 179121 164051
rect 179149 164023 194419 164051
rect 194447 164023 194481 164051
rect 194509 164023 209779 164051
rect 209807 164023 209841 164051
rect 209869 164023 225139 164051
rect 225167 164023 225201 164051
rect 225229 164023 240499 164051
rect 240527 164023 240561 164051
rect 240589 164023 255859 164051
rect 255887 164023 255921 164051
rect 255949 164023 271219 164051
rect 271247 164023 271281 164051
rect 271309 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298990 164051
rect -958 163989 298990 164023
rect -958 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 102259 163989
rect 102287 163961 102321 163989
rect 102349 163961 117619 163989
rect 117647 163961 117681 163989
rect 117709 163961 132979 163989
rect 133007 163961 133041 163989
rect 133069 163961 148339 163989
rect 148367 163961 148401 163989
rect 148429 163961 163699 163989
rect 163727 163961 163761 163989
rect 163789 163961 179059 163989
rect 179087 163961 179121 163989
rect 179149 163961 194419 163989
rect 194447 163961 194481 163989
rect 194509 163961 209779 163989
rect 209807 163961 209841 163989
rect 209869 163961 225139 163989
rect 225167 163961 225201 163989
rect 225229 163961 240499 163989
rect 240527 163961 240561 163989
rect 240589 163961 255859 163989
rect 255887 163961 255921 163989
rect 255949 163961 271219 163989
rect 271247 163961 271281 163989
rect 271309 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298990 163989
rect -958 163913 298990 163961
rect -958 158175 298990 158223
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 109939 158175
rect 109967 158147 110001 158175
rect 110029 158147 125299 158175
rect 125327 158147 125361 158175
rect 125389 158147 140659 158175
rect 140687 158147 140721 158175
rect 140749 158147 156019 158175
rect 156047 158147 156081 158175
rect 156109 158147 171379 158175
rect 171407 158147 171441 158175
rect 171469 158147 186739 158175
rect 186767 158147 186801 158175
rect 186829 158147 202099 158175
rect 202127 158147 202161 158175
rect 202189 158147 217459 158175
rect 217487 158147 217521 158175
rect 217549 158147 232819 158175
rect 232847 158147 232881 158175
rect 232909 158147 248179 158175
rect 248207 158147 248241 158175
rect 248269 158147 263539 158175
rect 263567 158147 263601 158175
rect 263629 158147 278899 158175
rect 278927 158147 278961 158175
rect 278989 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect -958 158113 298990 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 109939 158113
rect 109967 158085 110001 158113
rect 110029 158085 125299 158113
rect 125327 158085 125361 158113
rect 125389 158085 140659 158113
rect 140687 158085 140721 158113
rect 140749 158085 156019 158113
rect 156047 158085 156081 158113
rect 156109 158085 171379 158113
rect 171407 158085 171441 158113
rect 171469 158085 186739 158113
rect 186767 158085 186801 158113
rect 186829 158085 202099 158113
rect 202127 158085 202161 158113
rect 202189 158085 217459 158113
rect 217487 158085 217521 158113
rect 217549 158085 232819 158113
rect 232847 158085 232881 158113
rect 232909 158085 248179 158113
rect 248207 158085 248241 158113
rect 248269 158085 263539 158113
rect 263567 158085 263601 158113
rect 263629 158085 278899 158113
rect 278927 158085 278961 158113
rect 278989 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect -958 158051 298990 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 109939 158051
rect 109967 158023 110001 158051
rect 110029 158023 125299 158051
rect 125327 158023 125361 158051
rect 125389 158023 140659 158051
rect 140687 158023 140721 158051
rect 140749 158023 156019 158051
rect 156047 158023 156081 158051
rect 156109 158023 171379 158051
rect 171407 158023 171441 158051
rect 171469 158023 186739 158051
rect 186767 158023 186801 158051
rect 186829 158023 202099 158051
rect 202127 158023 202161 158051
rect 202189 158023 217459 158051
rect 217487 158023 217521 158051
rect 217549 158023 232819 158051
rect 232847 158023 232881 158051
rect 232909 158023 248179 158051
rect 248207 158023 248241 158051
rect 248269 158023 263539 158051
rect 263567 158023 263601 158051
rect 263629 158023 278899 158051
rect 278927 158023 278961 158051
rect 278989 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect -958 157989 298990 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 109939 157989
rect 109967 157961 110001 157989
rect 110029 157961 125299 157989
rect 125327 157961 125361 157989
rect 125389 157961 140659 157989
rect 140687 157961 140721 157989
rect 140749 157961 156019 157989
rect 156047 157961 156081 157989
rect 156109 157961 171379 157989
rect 171407 157961 171441 157989
rect 171469 157961 186739 157989
rect 186767 157961 186801 157989
rect 186829 157961 202099 157989
rect 202127 157961 202161 157989
rect 202189 157961 217459 157989
rect 217487 157961 217521 157989
rect 217549 157961 232819 157989
rect 232847 157961 232881 157989
rect 232909 157961 248179 157989
rect 248207 157961 248241 157989
rect 248269 157961 263539 157989
rect 263567 157961 263601 157989
rect 263629 157961 278899 157989
rect 278927 157961 278961 157989
rect 278989 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect -958 157913 298990 157961
rect -958 155175 298990 155223
rect -958 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 102259 155175
rect 102287 155147 102321 155175
rect 102349 155147 117619 155175
rect 117647 155147 117681 155175
rect 117709 155147 132979 155175
rect 133007 155147 133041 155175
rect 133069 155147 148339 155175
rect 148367 155147 148401 155175
rect 148429 155147 163699 155175
rect 163727 155147 163761 155175
rect 163789 155147 179059 155175
rect 179087 155147 179121 155175
rect 179149 155147 194419 155175
rect 194447 155147 194481 155175
rect 194509 155147 209779 155175
rect 209807 155147 209841 155175
rect 209869 155147 225139 155175
rect 225167 155147 225201 155175
rect 225229 155147 240499 155175
rect 240527 155147 240561 155175
rect 240589 155147 255859 155175
rect 255887 155147 255921 155175
rect 255949 155147 271219 155175
rect 271247 155147 271281 155175
rect 271309 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298990 155175
rect -958 155113 298990 155147
rect -958 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 102259 155113
rect 102287 155085 102321 155113
rect 102349 155085 117619 155113
rect 117647 155085 117681 155113
rect 117709 155085 132979 155113
rect 133007 155085 133041 155113
rect 133069 155085 148339 155113
rect 148367 155085 148401 155113
rect 148429 155085 163699 155113
rect 163727 155085 163761 155113
rect 163789 155085 179059 155113
rect 179087 155085 179121 155113
rect 179149 155085 194419 155113
rect 194447 155085 194481 155113
rect 194509 155085 209779 155113
rect 209807 155085 209841 155113
rect 209869 155085 225139 155113
rect 225167 155085 225201 155113
rect 225229 155085 240499 155113
rect 240527 155085 240561 155113
rect 240589 155085 255859 155113
rect 255887 155085 255921 155113
rect 255949 155085 271219 155113
rect 271247 155085 271281 155113
rect 271309 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298990 155113
rect -958 155051 298990 155085
rect -958 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 102259 155051
rect 102287 155023 102321 155051
rect 102349 155023 117619 155051
rect 117647 155023 117681 155051
rect 117709 155023 132979 155051
rect 133007 155023 133041 155051
rect 133069 155023 148339 155051
rect 148367 155023 148401 155051
rect 148429 155023 163699 155051
rect 163727 155023 163761 155051
rect 163789 155023 179059 155051
rect 179087 155023 179121 155051
rect 179149 155023 194419 155051
rect 194447 155023 194481 155051
rect 194509 155023 209779 155051
rect 209807 155023 209841 155051
rect 209869 155023 225139 155051
rect 225167 155023 225201 155051
rect 225229 155023 240499 155051
rect 240527 155023 240561 155051
rect 240589 155023 255859 155051
rect 255887 155023 255921 155051
rect 255949 155023 271219 155051
rect 271247 155023 271281 155051
rect 271309 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298990 155051
rect -958 154989 298990 155023
rect -958 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 102259 154989
rect 102287 154961 102321 154989
rect 102349 154961 117619 154989
rect 117647 154961 117681 154989
rect 117709 154961 132979 154989
rect 133007 154961 133041 154989
rect 133069 154961 148339 154989
rect 148367 154961 148401 154989
rect 148429 154961 163699 154989
rect 163727 154961 163761 154989
rect 163789 154961 179059 154989
rect 179087 154961 179121 154989
rect 179149 154961 194419 154989
rect 194447 154961 194481 154989
rect 194509 154961 209779 154989
rect 209807 154961 209841 154989
rect 209869 154961 225139 154989
rect 225167 154961 225201 154989
rect 225229 154961 240499 154989
rect 240527 154961 240561 154989
rect 240589 154961 255859 154989
rect 255887 154961 255921 154989
rect 255949 154961 271219 154989
rect 271247 154961 271281 154989
rect 271309 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298990 154989
rect -958 154913 298990 154961
rect -958 149175 298990 149223
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 109939 149175
rect 109967 149147 110001 149175
rect 110029 149147 125299 149175
rect 125327 149147 125361 149175
rect 125389 149147 140659 149175
rect 140687 149147 140721 149175
rect 140749 149147 156019 149175
rect 156047 149147 156081 149175
rect 156109 149147 171379 149175
rect 171407 149147 171441 149175
rect 171469 149147 186739 149175
rect 186767 149147 186801 149175
rect 186829 149147 202099 149175
rect 202127 149147 202161 149175
rect 202189 149147 217459 149175
rect 217487 149147 217521 149175
rect 217549 149147 232819 149175
rect 232847 149147 232881 149175
rect 232909 149147 248179 149175
rect 248207 149147 248241 149175
rect 248269 149147 263539 149175
rect 263567 149147 263601 149175
rect 263629 149147 278899 149175
rect 278927 149147 278961 149175
rect 278989 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect -958 149113 298990 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 109939 149113
rect 109967 149085 110001 149113
rect 110029 149085 125299 149113
rect 125327 149085 125361 149113
rect 125389 149085 140659 149113
rect 140687 149085 140721 149113
rect 140749 149085 156019 149113
rect 156047 149085 156081 149113
rect 156109 149085 171379 149113
rect 171407 149085 171441 149113
rect 171469 149085 186739 149113
rect 186767 149085 186801 149113
rect 186829 149085 202099 149113
rect 202127 149085 202161 149113
rect 202189 149085 217459 149113
rect 217487 149085 217521 149113
rect 217549 149085 232819 149113
rect 232847 149085 232881 149113
rect 232909 149085 248179 149113
rect 248207 149085 248241 149113
rect 248269 149085 263539 149113
rect 263567 149085 263601 149113
rect 263629 149085 278899 149113
rect 278927 149085 278961 149113
rect 278989 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect -958 149051 298990 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 109939 149051
rect 109967 149023 110001 149051
rect 110029 149023 125299 149051
rect 125327 149023 125361 149051
rect 125389 149023 140659 149051
rect 140687 149023 140721 149051
rect 140749 149023 156019 149051
rect 156047 149023 156081 149051
rect 156109 149023 171379 149051
rect 171407 149023 171441 149051
rect 171469 149023 186739 149051
rect 186767 149023 186801 149051
rect 186829 149023 202099 149051
rect 202127 149023 202161 149051
rect 202189 149023 217459 149051
rect 217487 149023 217521 149051
rect 217549 149023 232819 149051
rect 232847 149023 232881 149051
rect 232909 149023 248179 149051
rect 248207 149023 248241 149051
rect 248269 149023 263539 149051
rect 263567 149023 263601 149051
rect 263629 149023 278899 149051
rect 278927 149023 278961 149051
rect 278989 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect -958 148989 298990 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 109939 148989
rect 109967 148961 110001 148989
rect 110029 148961 125299 148989
rect 125327 148961 125361 148989
rect 125389 148961 140659 148989
rect 140687 148961 140721 148989
rect 140749 148961 156019 148989
rect 156047 148961 156081 148989
rect 156109 148961 171379 148989
rect 171407 148961 171441 148989
rect 171469 148961 186739 148989
rect 186767 148961 186801 148989
rect 186829 148961 202099 148989
rect 202127 148961 202161 148989
rect 202189 148961 217459 148989
rect 217487 148961 217521 148989
rect 217549 148961 232819 148989
rect 232847 148961 232881 148989
rect 232909 148961 248179 148989
rect 248207 148961 248241 148989
rect 248269 148961 263539 148989
rect 263567 148961 263601 148989
rect 263629 148961 278899 148989
rect 278927 148961 278961 148989
rect 278989 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect -958 148913 298990 148961
rect -958 146175 298990 146223
rect -958 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 102259 146175
rect 102287 146147 102321 146175
rect 102349 146147 117619 146175
rect 117647 146147 117681 146175
rect 117709 146147 132979 146175
rect 133007 146147 133041 146175
rect 133069 146147 148339 146175
rect 148367 146147 148401 146175
rect 148429 146147 163699 146175
rect 163727 146147 163761 146175
rect 163789 146147 179059 146175
rect 179087 146147 179121 146175
rect 179149 146147 194419 146175
rect 194447 146147 194481 146175
rect 194509 146147 209779 146175
rect 209807 146147 209841 146175
rect 209869 146147 225139 146175
rect 225167 146147 225201 146175
rect 225229 146147 240499 146175
rect 240527 146147 240561 146175
rect 240589 146147 255859 146175
rect 255887 146147 255921 146175
rect 255949 146147 271219 146175
rect 271247 146147 271281 146175
rect 271309 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298990 146175
rect -958 146113 298990 146147
rect -958 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 102259 146113
rect 102287 146085 102321 146113
rect 102349 146085 117619 146113
rect 117647 146085 117681 146113
rect 117709 146085 132979 146113
rect 133007 146085 133041 146113
rect 133069 146085 148339 146113
rect 148367 146085 148401 146113
rect 148429 146085 163699 146113
rect 163727 146085 163761 146113
rect 163789 146085 179059 146113
rect 179087 146085 179121 146113
rect 179149 146085 194419 146113
rect 194447 146085 194481 146113
rect 194509 146085 209779 146113
rect 209807 146085 209841 146113
rect 209869 146085 225139 146113
rect 225167 146085 225201 146113
rect 225229 146085 240499 146113
rect 240527 146085 240561 146113
rect 240589 146085 255859 146113
rect 255887 146085 255921 146113
rect 255949 146085 271219 146113
rect 271247 146085 271281 146113
rect 271309 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298990 146113
rect -958 146051 298990 146085
rect -958 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 102259 146051
rect 102287 146023 102321 146051
rect 102349 146023 117619 146051
rect 117647 146023 117681 146051
rect 117709 146023 132979 146051
rect 133007 146023 133041 146051
rect 133069 146023 148339 146051
rect 148367 146023 148401 146051
rect 148429 146023 163699 146051
rect 163727 146023 163761 146051
rect 163789 146023 179059 146051
rect 179087 146023 179121 146051
rect 179149 146023 194419 146051
rect 194447 146023 194481 146051
rect 194509 146023 209779 146051
rect 209807 146023 209841 146051
rect 209869 146023 225139 146051
rect 225167 146023 225201 146051
rect 225229 146023 240499 146051
rect 240527 146023 240561 146051
rect 240589 146023 255859 146051
rect 255887 146023 255921 146051
rect 255949 146023 271219 146051
rect 271247 146023 271281 146051
rect 271309 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298990 146051
rect -958 145989 298990 146023
rect -958 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 102259 145989
rect 102287 145961 102321 145989
rect 102349 145961 117619 145989
rect 117647 145961 117681 145989
rect 117709 145961 132979 145989
rect 133007 145961 133041 145989
rect 133069 145961 148339 145989
rect 148367 145961 148401 145989
rect 148429 145961 163699 145989
rect 163727 145961 163761 145989
rect 163789 145961 179059 145989
rect 179087 145961 179121 145989
rect 179149 145961 194419 145989
rect 194447 145961 194481 145989
rect 194509 145961 209779 145989
rect 209807 145961 209841 145989
rect 209869 145961 225139 145989
rect 225167 145961 225201 145989
rect 225229 145961 240499 145989
rect 240527 145961 240561 145989
rect 240589 145961 255859 145989
rect 255887 145961 255921 145989
rect 255949 145961 271219 145989
rect 271247 145961 271281 145989
rect 271309 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298990 145989
rect -958 145913 298990 145961
rect -958 140175 298990 140223
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 109939 140175
rect 109967 140147 110001 140175
rect 110029 140147 125299 140175
rect 125327 140147 125361 140175
rect 125389 140147 140659 140175
rect 140687 140147 140721 140175
rect 140749 140147 156019 140175
rect 156047 140147 156081 140175
rect 156109 140147 171379 140175
rect 171407 140147 171441 140175
rect 171469 140147 186739 140175
rect 186767 140147 186801 140175
rect 186829 140147 202099 140175
rect 202127 140147 202161 140175
rect 202189 140147 217459 140175
rect 217487 140147 217521 140175
rect 217549 140147 232819 140175
rect 232847 140147 232881 140175
rect 232909 140147 248179 140175
rect 248207 140147 248241 140175
rect 248269 140147 263539 140175
rect 263567 140147 263601 140175
rect 263629 140147 278899 140175
rect 278927 140147 278961 140175
rect 278989 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect -958 140113 298990 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 109939 140113
rect 109967 140085 110001 140113
rect 110029 140085 125299 140113
rect 125327 140085 125361 140113
rect 125389 140085 140659 140113
rect 140687 140085 140721 140113
rect 140749 140085 156019 140113
rect 156047 140085 156081 140113
rect 156109 140085 171379 140113
rect 171407 140085 171441 140113
rect 171469 140085 186739 140113
rect 186767 140085 186801 140113
rect 186829 140085 202099 140113
rect 202127 140085 202161 140113
rect 202189 140085 217459 140113
rect 217487 140085 217521 140113
rect 217549 140085 232819 140113
rect 232847 140085 232881 140113
rect 232909 140085 248179 140113
rect 248207 140085 248241 140113
rect 248269 140085 263539 140113
rect 263567 140085 263601 140113
rect 263629 140085 278899 140113
rect 278927 140085 278961 140113
rect 278989 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect -958 140051 298990 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 109939 140051
rect 109967 140023 110001 140051
rect 110029 140023 125299 140051
rect 125327 140023 125361 140051
rect 125389 140023 140659 140051
rect 140687 140023 140721 140051
rect 140749 140023 156019 140051
rect 156047 140023 156081 140051
rect 156109 140023 171379 140051
rect 171407 140023 171441 140051
rect 171469 140023 186739 140051
rect 186767 140023 186801 140051
rect 186829 140023 202099 140051
rect 202127 140023 202161 140051
rect 202189 140023 217459 140051
rect 217487 140023 217521 140051
rect 217549 140023 232819 140051
rect 232847 140023 232881 140051
rect 232909 140023 248179 140051
rect 248207 140023 248241 140051
rect 248269 140023 263539 140051
rect 263567 140023 263601 140051
rect 263629 140023 278899 140051
rect 278927 140023 278961 140051
rect 278989 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect -958 139989 298990 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 109939 139989
rect 109967 139961 110001 139989
rect 110029 139961 125299 139989
rect 125327 139961 125361 139989
rect 125389 139961 140659 139989
rect 140687 139961 140721 139989
rect 140749 139961 156019 139989
rect 156047 139961 156081 139989
rect 156109 139961 171379 139989
rect 171407 139961 171441 139989
rect 171469 139961 186739 139989
rect 186767 139961 186801 139989
rect 186829 139961 202099 139989
rect 202127 139961 202161 139989
rect 202189 139961 217459 139989
rect 217487 139961 217521 139989
rect 217549 139961 232819 139989
rect 232847 139961 232881 139989
rect 232909 139961 248179 139989
rect 248207 139961 248241 139989
rect 248269 139961 263539 139989
rect 263567 139961 263601 139989
rect 263629 139961 278899 139989
rect 278927 139961 278961 139989
rect 278989 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect -958 139913 298990 139961
rect -958 137175 298990 137223
rect -958 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 102259 137175
rect 102287 137147 102321 137175
rect 102349 137147 117619 137175
rect 117647 137147 117681 137175
rect 117709 137147 132979 137175
rect 133007 137147 133041 137175
rect 133069 137147 148339 137175
rect 148367 137147 148401 137175
rect 148429 137147 163699 137175
rect 163727 137147 163761 137175
rect 163789 137147 179059 137175
rect 179087 137147 179121 137175
rect 179149 137147 194419 137175
rect 194447 137147 194481 137175
rect 194509 137147 209779 137175
rect 209807 137147 209841 137175
rect 209869 137147 225139 137175
rect 225167 137147 225201 137175
rect 225229 137147 240499 137175
rect 240527 137147 240561 137175
rect 240589 137147 255859 137175
rect 255887 137147 255921 137175
rect 255949 137147 271219 137175
rect 271247 137147 271281 137175
rect 271309 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298990 137175
rect -958 137113 298990 137147
rect -958 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 102259 137113
rect 102287 137085 102321 137113
rect 102349 137085 117619 137113
rect 117647 137085 117681 137113
rect 117709 137085 132979 137113
rect 133007 137085 133041 137113
rect 133069 137085 148339 137113
rect 148367 137085 148401 137113
rect 148429 137085 163699 137113
rect 163727 137085 163761 137113
rect 163789 137085 179059 137113
rect 179087 137085 179121 137113
rect 179149 137085 194419 137113
rect 194447 137085 194481 137113
rect 194509 137085 209779 137113
rect 209807 137085 209841 137113
rect 209869 137085 225139 137113
rect 225167 137085 225201 137113
rect 225229 137085 240499 137113
rect 240527 137085 240561 137113
rect 240589 137085 255859 137113
rect 255887 137085 255921 137113
rect 255949 137085 271219 137113
rect 271247 137085 271281 137113
rect 271309 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298990 137113
rect -958 137051 298990 137085
rect -958 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 102259 137051
rect 102287 137023 102321 137051
rect 102349 137023 117619 137051
rect 117647 137023 117681 137051
rect 117709 137023 132979 137051
rect 133007 137023 133041 137051
rect 133069 137023 148339 137051
rect 148367 137023 148401 137051
rect 148429 137023 163699 137051
rect 163727 137023 163761 137051
rect 163789 137023 179059 137051
rect 179087 137023 179121 137051
rect 179149 137023 194419 137051
rect 194447 137023 194481 137051
rect 194509 137023 209779 137051
rect 209807 137023 209841 137051
rect 209869 137023 225139 137051
rect 225167 137023 225201 137051
rect 225229 137023 240499 137051
rect 240527 137023 240561 137051
rect 240589 137023 255859 137051
rect 255887 137023 255921 137051
rect 255949 137023 271219 137051
rect 271247 137023 271281 137051
rect 271309 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298990 137051
rect -958 136989 298990 137023
rect -958 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 102259 136989
rect 102287 136961 102321 136989
rect 102349 136961 117619 136989
rect 117647 136961 117681 136989
rect 117709 136961 132979 136989
rect 133007 136961 133041 136989
rect 133069 136961 148339 136989
rect 148367 136961 148401 136989
rect 148429 136961 163699 136989
rect 163727 136961 163761 136989
rect 163789 136961 179059 136989
rect 179087 136961 179121 136989
rect 179149 136961 194419 136989
rect 194447 136961 194481 136989
rect 194509 136961 209779 136989
rect 209807 136961 209841 136989
rect 209869 136961 225139 136989
rect 225167 136961 225201 136989
rect 225229 136961 240499 136989
rect 240527 136961 240561 136989
rect 240589 136961 255859 136989
rect 255887 136961 255921 136989
rect 255949 136961 271219 136989
rect 271247 136961 271281 136989
rect 271309 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298990 136989
rect -958 136913 298990 136961
rect -958 131175 298990 131223
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 109939 131175
rect 109967 131147 110001 131175
rect 110029 131147 125299 131175
rect 125327 131147 125361 131175
rect 125389 131147 140659 131175
rect 140687 131147 140721 131175
rect 140749 131147 156019 131175
rect 156047 131147 156081 131175
rect 156109 131147 171379 131175
rect 171407 131147 171441 131175
rect 171469 131147 186739 131175
rect 186767 131147 186801 131175
rect 186829 131147 202099 131175
rect 202127 131147 202161 131175
rect 202189 131147 217459 131175
rect 217487 131147 217521 131175
rect 217549 131147 232819 131175
rect 232847 131147 232881 131175
rect 232909 131147 248179 131175
rect 248207 131147 248241 131175
rect 248269 131147 263539 131175
rect 263567 131147 263601 131175
rect 263629 131147 278899 131175
rect 278927 131147 278961 131175
rect 278989 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect -958 131113 298990 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 109939 131113
rect 109967 131085 110001 131113
rect 110029 131085 125299 131113
rect 125327 131085 125361 131113
rect 125389 131085 140659 131113
rect 140687 131085 140721 131113
rect 140749 131085 156019 131113
rect 156047 131085 156081 131113
rect 156109 131085 171379 131113
rect 171407 131085 171441 131113
rect 171469 131085 186739 131113
rect 186767 131085 186801 131113
rect 186829 131085 202099 131113
rect 202127 131085 202161 131113
rect 202189 131085 217459 131113
rect 217487 131085 217521 131113
rect 217549 131085 232819 131113
rect 232847 131085 232881 131113
rect 232909 131085 248179 131113
rect 248207 131085 248241 131113
rect 248269 131085 263539 131113
rect 263567 131085 263601 131113
rect 263629 131085 278899 131113
rect 278927 131085 278961 131113
rect 278989 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect -958 131051 298990 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 109939 131051
rect 109967 131023 110001 131051
rect 110029 131023 125299 131051
rect 125327 131023 125361 131051
rect 125389 131023 140659 131051
rect 140687 131023 140721 131051
rect 140749 131023 156019 131051
rect 156047 131023 156081 131051
rect 156109 131023 171379 131051
rect 171407 131023 171441 131051
rect 171469 131023 186739 131051
rect 186767 131023 186801 131051
rect 186829 131023 202099 131051
rect 202127 131023 202161 131051
rect 202189 131023 217459 131051
rect 217487 131023 217521 131051
rect 217549 131023 232819 131051
rect 232847 131023 232881 131051
rect 232909 131023 248179 131051
rect 248207 131023 248241 131051
rect 248269 131023 263539 131051
rect 263567 131023 263601 131051
rect 263629 131023 278899 131051
rect 278927 131023 278961 131051
rect 278989 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect -958 130989 298990 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130961 109939 130989
rect 109967 130961 110001 130989
rect 110029 130961 125299 130989
rect 125327 130961 125361 130989
rect 125389 130961 140659 130989
rect 140687 130961 140721 130989
rect 140749 130961 156019 130989
rect 156047 130961 156081 130989
rect 156109 130961 171379 130989
rect 171407 130961 171441 130989
rect 171469 130961 186739 130989
rect 186767 130961 186801 130989
rect 186829 130961 202099 130989
rect 202127 130961 202161 130989
rect 202189 130961 217459 130989
rect 217487 130961 217521 130989
rect 217549 130961 232819 130989
rect 232847 130961 232881 130989
rect 232909 130961 248179 130989
rect 248207 130961 248241 130989
rect 248269 130961 263539 130989
rect 263567 130961 263601 130989
rect 263629 130961 278899 130989
rect 278927 130961 278961 130989
rect 278989 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect -958 130913 298990 130961
rect -958 128175 298990 128223
rect -958 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 102259 128175
rect 102287 128147 102321 128175
rect 102349 128147 117619 128175
rect 117647 128147 117681 128175
rect 117709 128147 132979 128175
rect 133007 128147 133041 128175
rect 133069 128147 148339 128175
rect 148367 128147 148401 128175
rect 148429 128147 163699 128175
rect 163727 128147 163761 128175
rect 163789 128147 179059 128175
rect 179087 128147 179121 128175
rect 179149 128147 194419 128175
rect 194447 128147 194481 128175
rect 194509 128147 209779 128175
rect 209807 128147 209841 128175
rect 209869 128147 225139 128175
rect 225167 128147 225201 128175
rect 225229 128147 240499 128175
rect 240527 128147 240561 128175
rect 240589 128147 255859 128175
rect 255887 128147 255921 128175
rect 255949 128147 271219 128175
rect 271247 128147 271281 128175
rect 271309 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298990 128175
rect -958 128113 298990 128147
rect -958 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 102259 128113
rect 102287 128085 102321 128113
rect 102349 128085 117619 128113
rect 117647 128085 117681 128113
rect 117709 128085 132979 128113
rect 133007 128085 133041 128113
rect 133069 128085 148339 128113
rect 148367 128085 148401 128113
rect 148429 128085 163699 128113
rect 163727 128085 163761 128113
rect 163789 128085 179059 128113
rect 179087 128085 179121 128113
rect 179149 128085 194419 128113
rect 194447 128085 194481 128113
rect 194509 128085 209779 128113
rect 209807 128085 209841 128113
rect 209869 128085 225139 128113
rect 225167 128085 225201 128113
rect 225229 128085 240499 128113
rect 240527 128085 240561 128113
rect 240589 128085 255859 128113
rect 255887 128085 255921 128113
rect 255949 128085 271219 128113
rect 271247 128085 271281 128113
rect 271309 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298990 128113
rect -958 128051 298990 128085
rect -958 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 102259 128051
rect 102287 128023 102321 128051
rect 102349 128023 117619 128051
rect 117647 128023 117681 128051
rect 117709 128023 132979 128051
rect 133007 128023 133041 128051
rect 133069 128023 148339 128051
rect 148367 128023 148401 128051
rect 148429 128023 163699 128051
rect 163727 128023 163761 128051
rect 163789 128023 179059 128051
rect 179087 128023 179121 128051
rect 179149 128023 194419 128051
rect 194447 128023 194481 128051
rect 194509 128023 209779 128051
rect 209807 128023 209841 128051
rect 209869 128023 225139 128051
rect 225167 128023 225201 128051
rect 225229 128023 240499 128051
rect 240527 128023 240561 128051
rect 240589 128023 255859 128051
rect 255887 128023 255921 128051
rect 255949 128023 271219 128051
rect 271247 128023 271281 128051
rect 271309 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298990 128051
rect -958 127989 298990 128023
rect -958 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 102259 127989
rect 102287 127961 102321 127989
rect 102349 127961 117619 127989
rect 117647 127961 117681 127989
rect 117709 127961 132979 127989
rect 133007 127961 133041 127989
rect 133069 127961 148339 127989
rect 148367 127961 148401 127989
rect 148429 127961 163699 127989
rect 163727 127961 163761 127989
rect 163789 127961 179059 127989
rect 179087 127961 179121 127989
rect 179149 127961 194419 127989
rect 194447 127961 194481 127989
rect 194509 127961 209779 127989
rect 209807 127961 209841 127989
rect 209869 127961 225139 127989
rect 225167 127961 225201 127989
rect 225229 127961 240499 127989
rect 240527 127961 240561 127989
rect 240589 127961 255859 127989
rect 255887 127961 255921 127989
rect 255949 127961 271219 127989
rect 271247 127961 271281 127989
rect 271309 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298990 127989
rect -958 127913 298990 127961
rect -958 122175 298990 122223
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 109939 122175
rect 109967 122147 110001 122175
rect 110029 122147 125299 122175
rect 125327 122147 125361 122175
rect 125389 122147 140659 122175
rect 140687 122147 140721 122175
rect 140749 122147 156019 122175
rect 156047 122147 156081 122175
rect 156109 122147 171379 122175
rect 171407 122147 171441 122175
rect 171469 122147 186739 122175
rect 186767 122147 186801 122175
rect 186829 122147 202099 122175
rect 202127 122147 202161 122175
rect 202189 122147 217459 122175
rect 217487 122147 217521 122175
rect 217549 122147 232819 122175
rect 232847 122147 232881 122175
rect 232909 122147 248179 122175
rect 248207 122147 248241 122175
rect 248269 122147 263539 122175
rect 263567 122147 263601 122175
rect 263629 122147 278899 122175
rect 278927 122147 278961 122175
rect 278989 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect -958 122113 298990 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 109939 122113
rect 109967 122085 110001 122113
rect 110029 122085 125299 122113
rect 125327 122085 125361 122113
rect 125389 122085 140659 122113
rect 140687 122085 140721 122113
rect 140749 122085 156019 122113
rect 156047 122085 156081 122113
rect 156109 122085 171379 122113
rect 171407 122085 171441 122113
rect 171469 122085 186739 122113
rect 186767 122085 186801 122113
rect 186829 122085 202099 122113
rect 202127 122085 202161 122113
rect 202189 122085 217459 122113
rect 217487 122085 217521 122113
rect 217549 122085 232819 122113
rect 232847 122085 232881 122113
rect 232909 122085 248179 122113
rect 248207 122085 248241 122113
rect 248269 122085 263539 122113
rect 263567 122085 263601 122113
rect 263629 122085 278899 122113
rect 278927 122085 278961 122113
rect 278989 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect -958 122051 298990 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 109939 122051
rect 109967 122023 110001 122051
rect 110029 122023 125299 122051
rect 125327 122023 125361 122051
rect 125389 122023 140659 122051
rect 140687 122023 140721 122051
rect 140749 122023 156019 122051
rect 156047 122023 156081 122051
rect 156109 122023 171379 122051
rect 171407 122023 171441 122051
rect 171469 122023 186739 122051
rect 186767 122023 186801 122051
rect 186829 122023 202099 122051
rect 202127 122023 202161 122051
rect 202189 122023 217459 122051
rect 217487 122023 217521 122051
rect 217549 122023 232819 122051
rect 232847 122023 232881 122051
rect 232909 122023 248179 122051
rect 248207 122023 248241 122051
rect 248269 122023 263539 122051
rect 263567 122023 263601 122051
rect 263629 122023 278899 122051
rect 278927 122023 278961 122051
rect 278989 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect -958 121989 298990 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 109939 121989
rect 109967 121961 110001 121989
rect 110029 121961 125299 121989
rect 125327 121961 125361 121989
rect 125389 121961 140659 121989
rect 140687 121961 140721 121989
rect 140749 121961 156019 121989
rect 156047 121961 156081 121989
rect 156109 121961 171379 121989
rect 171407 121961 171441 121989
rect 171469 121961 186739 121989
rect 186767 121961 186801 121989
rect 186829 121961 202099 121989
rect 202127 121961 202161 121989
rect 202189 121961 217459 121989
rect 217487 121961 217521 121989
rect 217549 121961 232819 121989
rect 232847 121961 232881 121989
rect 232909 121961 248179 121989
rect 248207 121961 248241 121989
rect 248269 121961 263539 121989
rect 263567 121961 263601 121989
rect 263629 121961 278899 121989
rect 278927 121961 278961 121989
rect 278989 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect -958 121913 298990 121961
rect -958 119175 298990 119223
rect -958 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 102259 119175
rect 102287 119147 102321 119175
rect 102349 119147 117619 119175
rect 117647 119147 117681 119175
rect 117709 119147 132979 119175
rect 133007 119147 133041 119175
rect 133069 119147 148339 119175
rect 148367 119147 148401 119175
rect 148429 119147 163699 119175
rect 163727 119147 163761 119175
rect 163789 119147 179059 119175
rect 179087 119147 179121 119175
rect 179149 119147 194419 119175
rect 194447 119147 194481 119175
rect 194509 119147 209779 119175
rect 209807 119147 209841 119175
rect 209869 119147 225139 119175
rect 225167 119147 225201 119175
rect 225229 119147 240499 119175
rect 240527 119147 240561 119175
rect 240589 119147 255859 119175
rect 255887 119147 255921 119175
rect 255949 119147 271219 119175
rect 271247 119147 271281 119175
rect 271309 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298990 119175
rect -958 119113 298990 119147
rect -958 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 102259 119113
rect 102287 119085 102321 119113
rect 102349 119085 117619 119113
rect 117647 119085 117681 119113
rect 117709 119085 132979 119113
rect 133007 119085 133041 119113
rect 133069 119085 148339 119113
rect 148367 119085 148401 119113
rect 148429 119085 163699 119113
rect 163727 119085 163761 119113
rect 163789 119085 179059 119113
rect 179087 119085 179121 119113
rect 179149 119085 194419 119113
rect 194447 119085 194481 119113
rect 194509 119085 209779 119113
rect 209807 119085 209841 119113
rect 209869 119085 225139 119113
rect 225167 119085 225201 119113
rect 225229 119085 240499 119113
rect 240527 119085 240561 119113
rect 240589 119085 255859 119113
rect 255887 119085 255921 119113
rect 255949 119085 271219 119113
rect 271247 119085 271281 119113
rect 271309 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298990 119113
rect -958 119051 298990 119085
rect -958 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 102259 119051
rect 102287 119023 102321 119051
rect 102349 119023 117619 119051
rect 117647 119023 117681 119051
rect 117709 119023 132979 119051
rect 133007 119023 133041 119051
rect 133069 119023 148339 119051
rect 148367 119023 148401 119051
rect 148429 119023 163699 119051
rect 163727 119023 163761 119051
rect 163789 119023 179059 119051
rect 179087 119023 179121 119051
rect 179149 119023 194419 119051
rect 194447 119023 194481 119051
rect 194509 119023 209779 119051
rect 209807 119023 209841 119051
rect 209869 119023 225139 119051
rect 225167 119023 225201 119051
rect 225229 119023 240499 119051
rect 240527 119023 240561 119051
rect 240589 119023 255859 119051
rect 255887 119023 255921 119051
rect 255949 119023 271219 119051
rect 271247 119023 271281 119051
rect 271309 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298990 119051
rect -958 118989 298990 119023
rect -958 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 102259 118989
rect 102287 118961 102321 118989
rect 102349 118961 117619 118989
rect 117647 118961 117681 118989
rect 117709 118961 132979 118989
rect 133007 118961 133041 118989
rect 133069 118961 148339 118989
rect 148367 118961 148401 118989
rect 148429 118961 163699 118989
rect 163727 118961 163761 118989
rect 163789 118961 179059 118989
rect 179087 118961 179121 118989
rect 179149 118961 194419 118989
rect 194447 118961 194481 118989
rect 194509 118961 209779 118989
rect 209807 118961 209841 118989
rect 209869 118961 225139 118989
rect 225167 118961 225201 118989
rect 225229 118961 240499 118989
rect 240527 118961 240561 118989
rect 240589 118961 255859 118989
rect 255887 118961 255921 118989
rect 255949 118961 271219 118989
rect 271247 118961 271281 118989
rect 271309 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298990 118989
rect -958 118913 298990 118961
rect -958 113175 298990 113223
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 109939 113175
rect 109967 113147 110001 113175
rect 110029 113147 125299 113175
rect 125327 113147 125361 113175
rect 125389 113147 140659 113175
rect 140687 113147 140721 113175
rect 140749 113147 156019 113175
rect 156047 113147 156081 113175
rect 156109 113147 171379 113175
rect 171407 113147 171441 113175
rect 171469 113147 186739 113175
rect 186767 113147 186801 113175
rect 186829 113147 202099 113175
rect 202127 113147 202161 113175
rect 202189 113147 217459 113175
rect 217487 113147 217521 113175
rect 217549 113147 232819 113175
rect 232847 113147 232881 113175
rect 232909 113147 248179 113175
rect 248207 113147 248241 113175
rect 248269 113147 263539 113175
rect 263567 113147 263601 113175
rect 263629 113147 278899 113175
rect 278927 113147 278961 113175
rect 278989 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect -958 113113 298990 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 109939 113113
rect 109967 113085 110001 113113
rect 110029 113085 125299 113113
rect 125327 113085 125361 113113
rect 125389 113085 140659 113113
rect 140687 113085 140721 113113
rect 140749 113085 156019 113113
rect 156047 113085 156081 113113
rect 156109 113085 171379 113113
rect 171407 113085 171441 113113
rect 171469 113085 186739 113113
rect 186767 113085 186801 113113
rect 186829 113085 202099 113113
rect 202127 113085 202161 113113
rect 202189 113085 217459 113113
rect 217487 113085 217521 113113
rect 217549 113085 232819 113113
rect 232847 113085 232881 113113
rect 232909 113085 248179 113113
rect 248207 113085 248241 113113
rect 248269 113085 263539 113113
rect 263567 113085 263601 113113
rect 263629 113085 278899 113113
rect 278927 113085 278961 113113
rect 278989 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect -958 113051 298990 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 109939 113051
rect 109967 113023 110001 113051
rect 110029 113023 125299 113051
rect 125327 113023 125361 113051
rect 125389 113023 140659 113051
rect 140687 113023 140721 113051
rect 140749 113023 156019 113051
rect 156047 113023 156081 113051
rect 156109 113023 171379 113051
rect 171407 113023 171441 113051
rect 171469 113023 186739 113051
rect 186767 113023 186801 113051
rect 186829 113023 202099 113051
rect 202127 113023 202161 113051
rect 202189 113023 217459 113051
rect 217487 113023 217521 113051
rect 217549 113023 232819 113051
rect 232847 113023 232881 113051
rect 232909 113023 248179 113051
rect 248207 113023 248241 113051
rect 248269 113023 263539 113051
rect 263567 113023 263601 113051
rect 263629 113023 278899 113051
rect 278927 113023 278961 113051
rect 278989 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect -958 112989 298990 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 109939 112989
rect 109967 112961 110001 112989
rect 110029 112961 125299 112989
rect 125327 112961 125361 112989
rect 125389 112961 140659 112989
rect 140687 112961 140721 112989
rect 140749 112961 156019 112989
rect 156047 112961 156081 112989
rect 156109 112961 171379 112989
rect 171407 112961 171441 112989
rect 171469 112961 186739 112989
rect 186767 112961 186801 112989
rect 186829 112961 202099 112989
rect 202127 112961 202161 112989
rect 202189 112961 217459 112989
rect 217487 112961 217521 112989
rect 217549 112961 232819 112989
rect 232847 112961 232881 112989
rect 232909 112961 248179 112989
rect 248207 112961 248241 112989
rect 248269 112961 263539 112989
rect 263567 112961 263601 112989
rect 263629 112961 278899 112989
rect 278927 112961 278961 112989
rect 278989 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect -958 112913 298990 112961
rect -958 110175 298990 110223
rect -958 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 102259 110175
rect 102287 110147 102321 110175
rect 102349 110147 117619 110175
rect 117647 110147 117681 110175
rect 117709 110147 132979 110175
rect 133007 110147 133041 110175
rect 133069 110147 148339 110175
rect 148367 110147 148401 110175
rect 148429 110147 163699 110175
rect 163727 110147 163761 110175
rect 163789 110147 179059 110175
rect 179087 110147 179121 110175
rect 179149 110147 194419 110175
rect 194447 110147 194481 110175
rect 194509 110147 209779 110175
rect 209807 110147 209841 110175
rect 209869 110147 225139 110175
rect 225167 110147 225201 110175
rect 225229 110147 240499 110175
rect 240527 110147 240561 110175
rect 240589 110147 255859 110175
rect 255887 110147 255921 110175
rect 255949 110147 271219 110175
rect 271247 110147 271281 110175
rect 271309 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298990 110175
rect -958 110113 298990 110147
rect -958 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 102259 110113
rect 102287 110085 102321 110113
rect 102349 110085 117619 110113
rect 117647 110085 117681 110113
rect 117709 110085 132979 110113
rect 133007 110085 133041 110113
rect 133069 110085 148339 110113
rect 148367 110085 148401 110113
rect 148429 110085 163699 110113
rect 163727 110085 163761 110113
rect 163789 110085 179059 110113
rect 179087 110085 179121 110113
rect 179149 110085 194419 110113
rect 194447 110085 194481 110113
rect 194509 110085 209779 110113
rect 209807 110085 209841 110113
rect 209869 110085 225139 110113
rect 225167 110085 225201 110113
rect 225229 110085 240499 110113
rect 240527 110085 240561 110113
rect 240589 110085 255859 110113
rect 255887 110085 255921 110113
rect 255949 110085 271219 110113
rect 271247 110085 271281 110113
rect 271309 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298990 110113
rect -958 110051 298990 110085
rect -958 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 102259 110051
rect 102287 110023 102321 110051
rect 102349 110023 117619 110051
rect 117647 110023 117681 110051
rect 117709 110023 132979 110051
rect 133007 110023 133041 110051
rect 133069 110023 148339 110051
rect 148367 110023 148401 110051
rect 148429 110023 163699 110051
rect 163727 110023 163761 110051
rect 163789 110023 179059 110051
rect 179087 110023 179121 110051
rect 179149 110023 194419 110051
rect 194447 110023 194481 110051
rect 194509 110023 209779 110051
rect 209807 110023 209841 110051
rect 209869 110023 225139 110051
rect 225167 110023 225201 110051
rect 225229 110023 240499 110051
rect 240527 110023 240561 110051
rect 240589 110023 255859 110051
rect 255887 110023 255921 110051
rect 255949 110023 271219 110051
rect 271247 110023 271281 110051
rect 271309 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298990 110051
rect -958 109989 298990 110023
rect -958 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 102259 109989
rect 102287 109961 102321 109989
rect 102349 109961 117619 109989
rect 117647 109961 117681 109989
rect 117709 109961 132979 109989
rect 133007 109961 133041 109989
rect 133069 109961 148339 109989
rect 148367 109961 148401 109989
rect 148429 109961 163699 109989
rect 163727 109961 163761 109989
rect 163789 109961 179059 109989
rect 179087 109961 179121 109989
rect 179149 109961 194419 109989
rect 194447 109961 194481 109989
rect 194509 109961 209779 109989
rect 209807 109961 209841 109989
rect 209869 109961 225139 109989
rect 225167 109961 225201 109989
rect 225229 109961 240499 109989
rect 240527 109961 240561 109989
rect 240589 109961 255859 109989
rect 255887 109961 255921 109989
rect 255949 109961 271219 109989
rect 271247 109961 271281 109989
rect 271309 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298990 109989
rect -958 109913 298990 109961
rect -958 104175 298990 104223
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 109939 104175
rect 109967 104147 110001 104175
rect 110029 104147 125299 104175
rect 125327 104147 125361 104175
rect 125389 104147 140659 104175
rect 140687 104147 140721 104175
rect 140749 104147 156019 104175
rect 156047 104147 156081 104175
rect 156109 104147 171379 104175
rect 171407 104147 171441 104175
rect 171469 104147 186739 104175
rect 186767 104147 186801 104175
rect 186829 104147 202099 104175
rect 202127 104147 202161 104175
rect 202189 104147 217459 104175
rect 217487 104147 217521 104175
rect 217549 104147 232819 104175
rect 232847 104147 232881 104175
rect 232909 104147 248179 104175
rect 248207 104147 248241 104175
rect 248269 104147 263539 104175
rect 263567 104147 263601 104175
rect 263629 104147 278899 104175
rect 278927 104147 278961 104175
rect 278989 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect -958 104113 298990 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 109939 104113
rect 109967 104085 110001 104113
rect 110029 104085 125299 104113
rect 125327 104085 125361 104113
rect 125389 104085 140659 104113
rect 140687 104085 140721 104113
rect 140749 104085 156019 104113
rect 156047 104085 156081 104113
rect 156109 104085 171379 104113
rect 171407 104085 171441 104113
rect 171469 104085 186739 104113
rect 186767 104085 186801 104113
rect 186829 104085 202099 104113
rect 202127 104085 202161 104113
rect 202189 104085 217459 104113
rect 217487 104085 217521 104113
rect 217549 104085 232819 104113
rect 232847 104085 232881 104113
rect 232909 104085 248179 104113
rect 248207 104085 248241 104113
rect 248269 104085 263539 104113
rect 263567 104085 263601 104113
rect 263629 104085 278899 104113
rect 278927 104085 278961 104113
rect 278989 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect -958 104051 298990 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 109939 104051
rect 109967 104023 110001 104051
rect 110029 104023 125299 104051
rect 125327 104023 125361 104051
rect 125389 104023 140659 104051
rect 140687 104023 140721 104051
rect 140749 104023 156019 104051
rect 156047 104023 156081 104051
rect 156109 104023 171379 104051
rect 171407 104023 171441 104051
rect 171469 104023 186739 104051
rect 186767 104023 186801 104051
rect 186829 104023 202099 104051
rect 202127 104023 202161 104051
rect 202189 104023 217459 104051
rect 217487 104023 217521 104051
rect 217549 104023 232819 104051
rect 232847 104023 232881 104051
rect 232909 104023 248179 104051
rect 248207 104023 248241 104051
rect 248269 104023 263539 104051
rect 263567 104023 263601 104051
rect 263629 104023 278899 104051
rect 278927 104023 278961 104051
rect 278989 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect -958 103989 298990 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 109939 103989
rect 109967 103961 110001 103989
rect 110029 103961 125299 103989
rect 125327 103961 125361 103989
rect 125389 103961 140659 103989
rect 140687 103961 140721 103989
rect 140749 103961 156019 103989
rect 156047 103961 156081 103989
rect 156109 103961 171379 103989
rect 171407 103961 171441 103989
rect 171469 103961 186739 103989
rect 186767 103961 186801 103989
rect 186829 103961 202099 103989
rect 202127 103961 202161 103989
rect 202189 103961 217459 103989
rect 217487 103961 217521 103989
rect 217549 103961 232819 103989
rect 232847 103961 232881 103989
rect 232909 103961 248179 103989
rect 248207 103961 248241 103989
rect 248269 103961 263539 103989
rect 263567 103961 263601 103989
rect 263629 103961 278899 103989
rect 278927 103961 278961 103989
rect 278989 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect -958 103913 298990 103961
rect -958 101175 298990 101223
rect -958 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298990 101175
rect -958 101113 298990 101147
rect -958 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298990 101113
rect -958 101051 298990 101085
rect -958 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298990 101051
rect -958 100989 298990 101023
rect -958 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298990 100989
rect -958 100913 298990 100961
rect -958 95175 298990 95223
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 173577 95175
rect 173605 95147 173639 95175
rect 173667 95147 173701 95175
rect 173729 95147 173763 95175
rect 173791 95147 188937 95175
rect 188965 95147 188999 95175
rect 189027 95147 189061 95175
rect 189089 95147 189123 95175
rect 189151 95147 204297 95175
rect 204325 95147 204359 95175
rect 204387 95147 204421 95175
rect 204449 95147 204483 95175
rect 204511 95147 219657 95175
rect 219685 95147 219719 95175
rect 219747 95147 219781 95175
rect 219809 95147 219843 95175
rect 219871 95147 235017 95175
rect 235045 95147 235079 95175
rect 235107 95147 235141 95175
rect 235169 95147 235203 95175
rect 235231 95147 250377 95175
rect 250405 95147 250439 95175
rect 250467 95147 250501 95175
rect 250529 95147 250563 95175
rect 250591 95147 265737 95175
rect 265765 95147 265799 95175
rect 265827 95147 265861 95175
rect 265889 95147 265923 95175
rect 265951 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect -958 95113 298990 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 173577 95113
rect 173605 95085 173639 95113
rect 173667 95085 173701 95113
rect 173729 95085 173763 95113
rect 173791 95085 188937 95113
rect 188965 95085 188999 95113
rect 189027 95085 189061 95113
rect 189089 95085 189123 95113
rect 189151 95085 204297 95113
rect 204325 95085 204359 95113
rect 204387 95085 204421 95113
rect 204449 95085 204483 95113
rect 204511 95085 219657 95113
rect 219685 95085 219719 95113
rect 219747 95085 219781 95113
rect 219809 95085 219843 95113
rect 219871 95085 235017 95113
rect 235045 95085 235079 95113
rect 235107 95085 235141 95113
rect 235169 95085 235203 95113
rect 235231 95085 250377 95113
rect 250405 95085 250439 95113
rect 250467 95085 250501 95113
rect 250529 95085 250563 95113
rect 250591 95085 265737 95113
rect 265765 95085 265799 95113
rect 265827 95085 265861 95113
rect 265889 95085 265923 95113
rect 265951 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect -958 95051 298990 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 173577 95051
rect 173605 95023 173639 95051
rect 173667 95023 173701 95051
rect 173729 95023 173763 95051
rect 173791 95023 188937 95051
rect 188965 95023 188999 95051
rect 189027 95023 189061 95051
rect 189089 95023 189123 95051
rect 189151 95023 204297 95051
rect 204325 95023 204359 95051
rect 204387 95023 204421 95051
rect 204449 95023 204483 95051
rect 204511 95023 219657 95051
rect 219685 95023 219719 95051
rect 219747 95023 219781 95051
rect 219809 95023 219843 95051
rect 219871 95023 235017 95051
rect 235045 95023 235079 95051
rect 235107 95023 235141 95051
rect 235169 95023 235203 95051
rect 235231 95023 250377 95051
rect 250405 95023 250439 95051
rect 250467 95023 250501 95051
rect 250529 95023 250563 95051
rect 250591 95023 265737 95051
rect 265765 95023 265799 95051
rect 265827 95023 265861 95051
rect 265889 95023 265923 95051
rect 265951 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect -958 94989 298990 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 173577 94989
rect 173605 94961 173639 94989
rect 173667 94961 173701 94989
rect 173729 94961 173763 94989
rect 173791 94961 188937 94989
rect 188965 94961 188999 94989
rect 189027 94961 189061 94989
rect 189089 94961 189123 94989
rect 189151 94961 204297 94989
rect 204325 94961 204359 94989
rect 204387 94961 204421 94989
rect 204449 94961 204483 94989
rect 204511 94961 219657 94989
rect 219685 94961 219719 94989
rect 219747 94961 219781 94989
rect 219809 94961 219843 94989
rect 219871 94961 235017 94989
rect 235045 94961 235079 94989
rect 235107 94961 235141 94989
rect 235169 94961 235203 94989
rect 235231 94961 250377 94989
rect 250405 94961 250439 94989
rect 250467 94961 250501 94989
rect 250529 94961 250563 94989
rect 250591 94961 265737 94989
rect 265765 94961 265799 94989
rect 265827 94961 265861 94989
rect 265889 94961 265923 94989
rect 265951 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect -958 94913 298990 94961
rect -958 92175 298990 92223
rect -958 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 171717 92175
rect 171745 92147 171779 92175
rect 171807 92147 171841 92175
rect 171869 92147 171903 92175
rect 171931 92147 187077 92175
rect 187105 92147 187139 92175
rect 187167 92147 187201 92175
rect 187229 92147 187263 92175
rect 187291 92147 202437 92175
rect 202465 92147 202499 92175
rect 202527 92147 202561 92175
rect 202589 92147 202623 92175
rect 202651 92147 217797 92175
rect 217825 92147 217859 92175
rect 217887 92147 217921 92175
rect 217949 92147 217983 92175
rect 218011 92147 233157 92175
rect 233185 92147 233219 92175
rect 233247 92147 233281 92175
rect 233309 92147 233343 92175
rect 233371 92147 248517 92175
rect 248545 92147 248579 92175
rect 248607 92147 248641 92175
rect 248669 92147 248703 92175
rect 248731 92147 263877 92175
rect 263905 92147 263939 92175
rect 263967 92147 264001 92175
rect 264029 92147 264063 92175
rect 264091 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298990 92175
rect -958 92113 298990 92147
rect -958 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 171717 92113
rect 171745 92085 171779 92113
rect 171807 92085 171841 92113
rect 171869 92085 171903 92113
rect 171931 92085 187077 92113
rect 187105 92085 187139 92113
rect 187167 92085 187201 92113
rect 187229 92085 187263 92113
rect 187291 92085 202437 92113
rect 202465 92085 202499 92113
rect 202527 92085 202561 92113
rect 202589 92085 202623 92113
rect 202651 92085 217797 92113
rect 217825 92085 217859 92113
rect 217887 92085 217921 92113
rect 217949 92085 217983 92113
rect 218011 92085 233157 92113
rect 233185 92085 233219 92113
rect 233247 92085 233281 92113
rect 233309 92085 233343 92113
rect 233371 92085 248517 92113
rect 248545 92085 248579 92113
rect 248607 92085 248641 92113
rect 248669 92085 248703 92113
rect 248731 92085 263877 92113
rect 263905 92085 263939 92113
rect 263967 92085 264001 92113
rect 264029 92085 264063 92113
rect 264091 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298990 92113
rect -958 92051 298990 92085
rect -958 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 171717 92051
rect 171745 92023 171779 92051
rect 171807 92023 171841 92051
rect 171869 92023 171903 92051
rect 171931 92023 187077 92051
rect 187105 92023 187139 92051
rect 187167 92023 187201 92051
rect 187229 92023 187263 92051
rect 187291 92023 202437 92051
rect 202465 92023 202499 92051
rect 202527 92023 202561 92051
rect 202589 92023 202623 92051
rect 202651 92023 217797 92051
rect 217825 92023 217859 92051
rect 217887 92023 217921 92051
rect 217949 92023 217983 92051
rect 218011 92023 233157 92051
rect 233185 92023 233219 92051
rect 233247 92023 233281 92051
rect 233309 92023 233343 92051
rect 233371 92023 248517 92051
rect 248545 92023 248579 92051
rect 248607 92023 248641 92051
rect 248669 92023 248703 92051
rect 248731 92023 263877 92051
rect 263905 92023 263939 92051
rect 263967 92023 264001 92051
rect 264029 92023 264063 92051
rect 264091 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298990 92051
rect -958 91989 298990 92023
rect -958 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 171717 91989
rect 171745 91961 171779 91989
rect 171807 91961 171841 91989
rect 171869 91961 171903 91989
rect 171931 91961 187077 91989
rect 187105 91961 187139 91989
rect 187167 91961 187201 91989
rect 187229 91961 187263 91989
rect 187291 91961 202437 91989
rect 202465 91961 202499 91989
rect 202527 91961 202561 91989
rect 202589 91961 202623 91989
rect 202651 91961 217797 91989
rect 217825 91961 217859 91989
rect 217887 91961 217921 91989
rect 217949 91961 217983 91989
rect 218011 91961 233157 91989
rect 233185 91961 233219 91989
rect 233247 91961 233281 91989
rect 233309 91961 233343 91989
rect 233371 91961 248517 91989
rect 248545 91961 248579 91989
rect 248607 91961 248641 91989
rect 248669 91961 248703 91989
rect 248731 91961 263877 91989
rect 263905 91961 263939 91989
rect 263967 91961 264001 91989
rect 264029 91961 264063 91989
rect 264091 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298990 91989
rect -958 91913 298990 91961
rect -958 86175 298990 86223
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 35337 86175
rect 35365 86147 35399 86175
rect 35427 86147 35461 86175
rect 35489 86147 35523 86175
rect 35551 86147 50697 86175
rect 50725 86147 50759 86175
rect 50787 86147 50821 86175
rect 50849 86147 50883 86175
rect 50911 86147 66057 86175
rect 66085 86147 66119 86175
rect 66147 86147 66181 86175
rect 66209 86147 66243 86175
rect 66271 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 173577 86175
rect 173605 86147 173639 86175
rect 173667 86147 173701 86175
rect 173729 86147 173763 86175
rect 173791 86147 188937 86175
rect 188965 86147 188999 86175
rect 189027 86147 189061 86175
rect 189089 86147 189123 86175
rect 189151 86147 204297 86175
rect 204325 86147 204359 86175
rect 204387 86147 204421 86175
rect 204449 86147 204483 86175
rect 204511 86147 219657 86175
rect 219685 86147 219719 86175
rect 219747 86147 219781 86175
rect 219809 86147 219843 86175
rect 219871 86147 235017 86175
rect 235045 86147 235079 86175
rect 235107 86147 235141 86175
rect 235169 86147 235203 86175
rect 235231 86147 250377 86175
rect 250405 86147 250439 86175
rect 250467 86147 250501 86175
rect 250529 86147 250563 86175
rect 250591 86147 265737 86175
rect 265765 86147 265799 86175
rect 265827 86147 265861 86175
rect 265889 86147 265923 86175
rect 265951 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect -958 86113 298990 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 35337 86113
rect 35365 86085 35399 86113
rect 35427 86085 35461 86113
rect 35489 86085 35523 86113
rect 35551 86085 50697 86113
rect 50725 86085 50759 86113
rect 50787 86085 50821 86113
rect 50849 86085 50883 86113
rect 50911 86085 66057 86113
rect 66085 86085 66119 86113
rect 66147 86085 66181 86113
rect 66209 86085 66243 86113
rect 66271 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 173577 86113
rect 173605 86085 173639 86113
rect 173667 86085 173701 86113
rect 173729 86085 173763 86113
rect 173791 86085 188937 86113
rect 188965 86085 188999 86113
rect 189027 86085 189061 86113
rect 189089 86085 189123 86113
rect 189151 86085 204297 86113
rect 204325 86085 204359 86113
rect 204387 86085 204421 86113
rect 204449 86085 204483 86113
rect 204511 86085 219657 86113
rect 219685 86085 219719 86113
rect 219747 86085 219781 86113
rect 219809 86085 219843 86113
rect 219871 86085 235017 86113
rect 235045 86085 235079 86113
rect 235107 86085 235141 86113
rect 235169 86085 235203 86113
rect 235231 86085 250377 86113
rect 250405 86085 250439 86113
rect 250467 86085 250501 86113
rect 250529 86085 250563 86113
rect 250591 86085 265737 86113
rect 265765 86085 265799 86113
rect 265827 86085 265861 86113
rect 265889 86085 265923 86113
rect 265951 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect -958 86051 298990 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 35337 86051
rect 35365 86023 35399 86051
rect 35427 86023 35461 86051
rect 35489 86023 35523 86051
rect 35551 86023 50697 86051
rect 50725 86023 50759 86051
rect 50787 86023 50821 86051
rect 50849 86023 50883 86051
rect 50911 86023 66057 86051
rect 66085 86023 66119 86051
rect 66147 86023 66181 86051
rect 66209 86023 66243 86051
rect 66271 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 173577 86051
rect 173605 86023 173639 86051
rect 173667 86023 173701 86051
rect 173729 86023 173763 86051
rect 173791 86023 188937 86051
rect 188965 86023 188999 86051
rect 189027 86023 189061 86051
rect 189089 86023 189123 86051
rect 189151 86023 204297 86051
rect 204325 86023 204359 86051
rect 204387 86023 204421 86051
rect 204449 86023 204483 86051
rect 204511 86023 219657 86051
rect 219685 86023 219719 86051
rect 219747 86023 219781 86051
rect 219809 86023 219843 86051
rect 219871 86023 235017 86051
rect 235045 86023 235079 86051
rect 235107 86023 235141 86051
rect 235169 86023 235203 86051
rect 235231 86023 250377 86051
rect 250405 86023 250439 86051
rect 250467 86023 250501 86051
rect 250529 86023 250563 86051
rect 250591 86023 265737 86051
rect 265765 86023 265799 86051
rect 265827 86023 265861 86051
rect 265889 86023 265923 86051
rect 265951 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect -958 85989 298990 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 35337 85989
rect 35365 85961 35399 85989
rect 35427 85961 35461 85989
rect 35489 85961 35523 85989
rect 35551 85961 50697 85989
rect 50725 85961 50759 85989
rect 50787 85961 50821 85989
rect 50849 85961 50883 85989
rect 50911 85961 66057 85989
rect 66085 85961 66119 85989
rect 66147 85961 66181 85989
rect 66209 85961 66243 85989
rect 66271 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 173577 85989
rect 173605 85961 173639 85989
rect 173667 85961 173701 85989
rect 173729 85961 173763 85989
rect 173791 85961 188937 85989
rect 188965 85961 188999 85989
rect 189027 85961 189061 85989
rect 189089 85961 189123 85989
rect 189151 85961 204297 85989
rect 204325 85961 204359 85989
rect 204387 85961 204421 85989
rect 204449 85961 204483 85989
rect 204511 85961 219657 85989
rect 219685 85961 219719 85989
rect 219747 85961 219781 85989
rect 219809 85961 219843 85989
rect 219871 85961 235017 85989
rect 235045 85961 235079 85989
rect 235107 85961 235141 85989
rect 235169 85961 235203 85989
rect 235231 85961 250377 85989
rect 250405 85961 250439 85989
rect 250467 85961 250501 85989
rect 250529 85961 250563 85989
rect 250591 85961 265737 85989
rect 265765 85961 265799 85989
rect 265827 85961 265861 85989
rect 265889 85961 265923 85989
rect 265951 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect -958 85913 298990 85961
rect -958 83175 298990 83223
rect -958 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 33477 83175
rect 33505 83147 33539 83175
rect 33567 83147 33601 83175
rect 33629 83147 33663 83175
rect 33691 83147 48837 83175
rect 48865 83147 48899 83175
rect 48927 83147 48961 83175
rect 48989 83147 49023 83175
rect 49051 83147 64197 83175
rect 64225 83147 64259 83175
rect 64287 83147 64321 83175
rect 64349 83147 64383 83175
rect 64411 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 171717 83175
rect 171745 83147 171779 83175
rect 171807 83147 171841 83175
rect 171869 83147 171903 83175
rect 171931 83147 187077 83175
rect 187105 83147 187139 83175
rect 187167 83147 187201 83175
rect 187229 83147 187263 83175
rect 187291 83147 202437 83175
rect 202465 83147 202499 83175
rect 202527 83147 202561 83175
rect 202589 83147 202623 83175
rect 202651 83147 217797 83175
rect 217825 83147 217859 83175
rect 217887 83147 217921 83175
rect 217949 83147 217983 83175
rect 218011 83147 233157 83175
rect 233185 83147 233219 83175
rect 233247 83147 233281 83175
rect 233309 83147 233343 83175
rect 233371 83147 248517 83175
rect 248545 83147 248579 83175
rect 248607 83147 248641 83175
rect 248669 83147 248703 83175
rect 248731 83147 263877 83175
rect 263905 83147 263939 83175
rect 263967 83147 264001 83175
rect 264029 83147 264063 83175
rect 264091 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298990 83175
rect -958 83113 298990 83147
rect -958 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 33477 83113
rect 33505 83085 33539 83113
rect 33567 83085 33601 83113
rect 33629 83085 33663 83113
rect 33691 83085 48837 83113
rect 48865 83085 48899 83113
rect 48927 83085 48961 83113
rect 48989 83085 49023 83113
rect 49051 83085 64197 83113
rect 64225 83085 64259 83113
rect 64287 83085 64321 83113
rect 64349 83085 64383 83113
rect 64411 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 171717 83113
rect 171745 83085 171779 83113
rect 171807 83085 171841 83113
rect 171869 83085 171903 83113
rect 171931 83085 187077 83113
rect 187105 83085 187139 83113
rect 187167 83085 187201 83113
rect 187229 83085 187263 83113
rect 187291 83085 202437 83113
rect 202465 83085 202499 83113
rect 202527 83085 202561 83113
rect 202589 83085 202623 83113
rect 202651 83085 217797 83113
rect 217825 83085 217859 83113
rect 217887 83085 217921 83113
rect 217949 83085 217983 83113
rect 218011 83085 233157 83113
rect 233185 83085 233219 83113
rect 233247 83085 233281 83113
rect 233309 83085 233343 83113
rect 233371 83085 248517 83113
rect 248545 83085 248579 83113
rect 248607 83085 248641 83113
rect 248669 83085 248703 83113
rect 248731 83085 263877 83113
rect 263905 83085 263939 83113
rect 263967 83085 264001 83113
rect 264029 83085 264063 83113
rect 264091 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298990 83113
rect -958 83051 298990 83085
rect -958 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 33477 83051
rect 33505 83023 33539 83051
rect 33567 83023 33601 83051
rect 33629 83023 33663 83051
rect 33691 83023 48837 83051
rect 48865 83023 48899 83051
rect 48927 83023 48961 83051
rect 48989 83023 49023 83051
rect 49051 83023 64197 83051
rect 64225 83023 64259 83051
rect 64287 83023 64321 83051
rect 64349 83023 64383 83051
rect 64411 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 171717 83051
rect 171745 83023 171779 83051
rect 171807 83023 171841 83051
rect 171869 83023 171903 83051
rect 171931 83023 187077 83051
rect 187105 83023 187139 83051
rect 187167 83023 187201 83051
rect 187229 83023 187263 83051
rect 187291 83023 202437 83051
rect 202465 83023 202499 83051
rect 202527 83023 202561 83051
rect 202589 83023 202623 83051
rect 202651 83023 217797 83051
rect 217825 83023 217859 83051
rect 217887 83023 217921 83051
rect 217949 83023 217983 83051
rect 218011 83023 233157 83051
rect 233185 83023 233219 83051
rect 233247 83023 233281 83051
rect 233309 83023 233343 83051
rect 233371 83023 248517 83051
rect 248545 83023 248579 83051
rect 248607 83023 248641 83051
rect 248669 83023 248703 83051
rect 248731 83023 263877 83051
rect 263905 83023 263939 83051
rect 263967 83023 264001 83051
rect 264029 83023 264063 83051
rect 264091 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298990 83051
rect -958 82989 298990 83023
rect -958 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 33477 82989
rect 33505 82961 33539 82989
rect 33567 82961 33601 82989
rect 33629 82961 33663 82989
rect 33691 82961 48837 82989
rect 48865 82961 48899 82989
rect 48927 82961 48961 82989
rect 48989 82961 49023 82989
rect 49051 82961 64197 82989
rect 64225 82961 64259 82989
rect 64287 82961 64321 82989
rect 64349 82961 64383 82989
rect 64411 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 171717 82989
rect 171745 82961 171779 82989
rect 171807 82961 171841 82989
rect 171869 82961 171903 82989
rect 171931 82961 187077 82989
rect 187105 82961 187139 82989
rect 187167 82961 187201 82989
rect 187229 82961 187263 82989
rect 187291 82961 202437 82989
rect 202465 82961 202499 82989
rect 202527 82961 202561 82989
rect 202589 82961 202623 82989
rect 202651 82961 217797 82989
rect 217825 82961 217859 82989
rect 217887 82961 217921 82989
rect 217949 82961 217983 82989
rect 218011 82961 233157 82989
rect 233185 82961 233219 82989
rect 233247 82961 233281 82989
rect 233309 82961 233343 82989
rect 233371 82961 248517 82989
rect 248545 82961 248579 82989
rect 248607 82961 248641 82989
rect 248669 82961 248703 82989
rect 248731 82961 263877 82989
rect 263905 82961 263939 82989
rect 263967 82961 264001 82989
rect 264029 82961 264063 82989
rect 264091 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298990 82989
rect -958 82913 298990 82961
rect -958 77175 298990 77223
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 35337 77175
rect 35365 77147 35399 77175
rect 35427 77147 35461 77175
rect 35489 77147 35523 77175
rect 35551 77147 50697 77175
rect 50725 77147 50759 77175
rect 50787 77147 50821 77175
rect 50849 77147 50883 77175
rect 50911 77147 66057 77175
rect 66085 77147 66119 77175
rect 66147 77147 66181 77175
rect 66209 77147 66243 77175
rect 66271 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 173577 77175
rect 173605 77147 173639 77175
rect 173667 77147 173701 77175
rect 173729 77147 173763 77175
rect 173791 77147 188937 77175
rect 188965 77147 188999 77175
rect 189027 77147 189061 77175
rect 189089 77147 189123 77175
rect 189151 77147 204297 77175
rect 204325 77147 204359 77175
rect 204387 77147 204421 77175
rect 204449 77147 204483 77175
rect 204511 77147 219657 77175
rect 219685 77147 219719 77175
rect 219747 77147 219781 77175
rect 219809 77147 219843 77175
rect 219871 77147 235017 77175
rect 235045 77147 235079 77175
rect 235107 77147 235141 77175
rect 235169 77147 235203 77175
rect 235231 77147 250377 77175
rect 250405 77147 250439 77175
rect 250467 77147 250501 77175
rect 250529 77147 250563 77175
rect 250591 77147 265737 77175
rect 265765 77147 265799 77175
rect 265827 77147 265861 77175
rect 265889 77147 265923 77175
rect 265951 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect -958 77113 298990 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 35337 77113
rect 35365 77085 35399 77113
rect 35427 77085 35461 77113
rect 35489 77085 35523 77113
rect 35551 77085 50697 77113
rect 50725 77085 50759 77113
rect 50787 77085 50821 77113
rect 50849 77085 50883 77113
rect 50911 77085 66057 77113
rect 66085 77085 66119 77113
rect 66147 77085 66181 77113
rect 66209 77085 66243 77113
rect 66271 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 173577 77113
rect 173605 77085 173639 77113
rect 173667 77085 173701 77113
rect 173729 77085 173763 77113
rect 173791 77085 188937 77113
rect 188965 77085 188999 77113
rect 189027 77085 189061 77113
rect 189089 77085 189123 77113
rect 189151 77085 204297 77113
rect 204325 77085 204359 77113
rect 204387 77085 204421 77113
rect 204449 77085 204483 77113
rect 204511 77085 219657 77113
rect 219685 77085 219719 77113
rect 219747 77085 219781 77113
rect 219809 77085 219843 77113
rect 219871 77085 235017 77113
rect 235045 77085 235079 77113
rect 235107 77085 235141 77113
rect 235169 77085 235203 77113
rect 235231 77085 250377 77113
rect 250405 77085 250439 77113
rect 250467 77085 250501 77113
rect 250529 77085 250563 77113
rect 250591 77085 265737 77113
rect 265765 77085 265799 77113
rect 265827 77085 265861 77113
rect 265889 77085 265923 77113
rect 265951 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect -958 77051 298990 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 35337 77051
rect 35365 77023 35399 77051
rect 35427 77023 35461 77051
rect 35489 77023 35523 77051
rect 35551 77023 50697 77051
rect 50725 77023 50759 77051
rect 50787 77023 50821 77051
rect 50849 77023 50883 77051
rect 50911 77023 66057 77051
rect 66085 77023 66119 77051
rect 66147 77023 66181 77051
rect 66209 77023 66243 77051
rect 66271 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 173577 77051
rect 173605 77023 173639 77051
rect 173667 77023 173701 77051
rect 173729 77023 173763 77051
rect 173791 77023 188937 77051
rect 188965 77023 188999 77051
rect 189027 77023 189061 77051
rect 189089 77023 189123 77051
rect 189151 77023 204297 77051
rect 204325 77023 204359 77051
rect 204387 77023 204421 77051
rect 204449 77023 204483 77051
rect 204511 77023 219657 77051
rect 219685 77023 219719 77051
rect 219747 77023 219781 77051
rect 219809 77023 219843 77051
rect 219871 77023 235017 77051
rect 235045 77023 235079 77051
rect 235107 77023 235141 77051
rect 235169 77023 235203 77051
rect 235231 77023 250377 77051
rect 250405 77023 250439 77051
rect 250467 77023 250501 77051
rect 250529 77023 250563 77051
rect 250591 77023 265737 77051
rect 265765 77023 265799 77051
rect 265827 77023 265861 77051
rect 265889 77023 265923 77051
rect 265951 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect -958 76989 298990 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 35337 76989
rect 35365 76961 35399 76989
rect 35427 76961 35461 76989
rect 35489 76961 35523 76989
rect 35551 76961 50697 76989
rect 50725 76961 50759 76989
rect 50787 76961 50821 76989
rect 50849 76961 50883 76989
rect 50911 76961 66057 76989
rect 66085 76961 66119 76989
rect 66147 76961 66181 76989
rect 66209 76961 66243 76989
rect 66271 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 173577 76989
rect 173605 76961 173639 76989
rect 173667 76961 173701 76989
rect 173729 76961 173763 76989
rect 173791 76961 188937 76989
rect 188965 76961 188999 76989
rect 189027 76961 189061 76989
rect 189089 76961 189123 76989
rect 189151 76961 204297 76989
rect 204325 76961 204359 76989
rect 204387 76961 204421 76989
rect 204449 76961 204483 76989
rect 204511 76961 219657 76989
rect 219685 76961 219719 76989
rect 219747 76961 219781 76989
rect 219809 76961 219843 76989
rect 219871 76961 235017 76989
rect 235045 76961 235079 76989
rect 235107 76961 235141 76989
rect 235169 76961 235203 76989
rect 235231 76961 250377 76989
rect 250405 76961 250439 76989
rect 250467 76961 250501 76989
rect 250529 76961 250563 76989
rect 250591 76961 265737 76989
rect 265765 76961 265799 76989
rect 265827 76961 265861 76989
rect 265889 76961 265923 76989
rect 265951 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect -958 76913 298990 76961
rect -958 74175 298990 74223
rect -958 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 171717 74175
rect 171745 74147 171779 74175
rect 171807 74147 171841 74175
rect 171869 74147 171903 74175
rect 171931 74147 187077 74175
rect 187105 74147 187139 74175
rect 187167 74147 187201 74175
rect 187229 74147 187263 74175
rect 187291 74147 202437 74175
rect 202465 74147 202499 74175
rect 202527 74147 202561 74175
rect 202589 74147 202623 74175
rect 202651 74147 217797 74175
rect 217825 74147 217859 74175
rect 217887 74147 217921 74175
rect 217949 74147 217983 74175
rect 218011 74147 233157 74175
rect 233185 74147 233219 74175
rect 233247 74147 233281 74175
rect 233309 74147 233343 74175
rect 233371 74147 248517 74175
rect 248545 74147 248579 74175
rect 248607 74147 248641 74175
rect 248669 74147 248703 74175
rect 248731 74147 263877 74175
rect 263905 74147 263939 74175
rect 263967 74147 264001 74175
rect 264029 74147 264063 74175
rect 264091 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298990 74175
rect -958 74113 298990 74147
rect -958 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 171717 74113
rect 171745 74085 171779 74113
rect 171807 74085 171841 74113
rect 171869 74085 171903 74113
rect 171931 74085 187077 74113
rect 187105 74085 187139 74113
rect 187167 74085 187201 74113
rect 187229 74085 187263 74113
rect 187291 74085 202437 74113
rect 202465 74085 202499 74113
rect 202527 74085 202561 74113
rect 202589 74085 202623 74113
rect 202651 74085 217797 74113
rect 217825 74085 217859 74113
rect 217887 74085 217921 74113
rect 217949 74085 217983 74113
rect 218011 74085 233157 74113
rect 233185 74085 233219 74113
rect 233247 74085 233281 74113
rect 233309 74085 233343 74113
rect 233371 74085 248517 74113
rect 248545 74085 248579 74113
rect 248607 74085 248641 74113
rect 248669 74085 248703 74113
rect 248731 74085 263877 74113
rect 263905 74085 263939 74113
rect 263967 74085 264001 74113
rect 264029 74085 264063 74113
rect 264091 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298990 74113
rect -958 74051 298990 74085
rect -958 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 171717 74051
rect 171745 74023 171779 74051
rect 171807 74023 171841 74051
rect 171869 74023 171903 74051
rect 171931 74023 187077 74051
rect 187105 74023 187139 74051
rect 187167 74023 187201 74051
rect 187229 74023 187263 74051
rect 187291 74023 202437 74051
rect 202465 74023 202499 74051
rect 202527 74023 202561 74051
rect 202589 74023 202623 74051
rect 202651 74023 217797 74051
rect 217825 74023 217859 74051
rect 217887 74023 217921 74051
rect 217949 74023 217983 74051
rect 218011 74023 233157 74051
rect 233185 74023 233219 74051
rect 233247 74023 233281 74051
rect 233309 74023 233343 74051
rect 233371 74023 248517 74051
rect 248545 74023 248579 74051
rect 248607 74023 248641 74051
rect 248669 74023 248703 74051
rect 248731 74023 263877 74051
rect 263905 74023 263939 74051
rect 263967 74023 264001 74051
rect 264029 74023 264063 74051
rect 264091 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298990 74051
rect -958 73989 298990 74023
rect -958 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 171717 73989
rect 171745 73961 171779 73989
rect 171807 73961 171841 73989
rect 171869 73961 171903 73989
rect 171931 73961 187077 73989
rect 187105 73961 187139 73989
rect 187167 73961 187201 73989
rect 187229 73961 187263 73989
rect 187291 73961 202437 73989
rect 202465 73961 202499 73989
rect 202527 73961 202561 73989
rect 202589 73961 202623 73989
rect 202651 73961 217797 73989
rect 217825 73961 217859 73989
rect 217887 73961 217921 73989
rect 217949 73961 217983 73989
rect 218011 73961 233157 73989
rect 233185 73961 233219 73989
rect 233247 73961 233281 73989
rect 233309 73961 233343 73989
rect 233371 73961 248517 73989
rect 248545 73961 248579 73989
rect 248607 73961 248641 73989
rect 248669 73961 248703 73989
rect 248731 73961 263877 73989
rect 263905 73961 263939 73989
rect 263967 73961 264001 73989
rect 264029 73961 264063 73989
rect 264091 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298990 73989
rect -958 73913 298990 73961
rect -958 68175 298990 68223
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 173577 68175
rect 173605 68147 173639 68175
rect 173667 68147 173701 68175
rect 173729 68147 173763 68175
rect 173791 68147 188937 68175
rect 188965 68147 188999 68175
rect 189027 68147 189061 68175
rect 189089 68147 189123 68175
rect 189151 68147 204297 68175
rect 204325 68147 204359 68175
rect 204387 68147 204421 68175
rect 204449 68147 204483 68175
rect 204511 68147 219657 68175
rect 219685 68147 219719 68175
rect 219747 68147 219781 68175
rect 219809 68147 219843 68175
rect 219871 68147 235017 68175
rect 235045 68147 235079 68175
rect 235107 68147 235141 68175
rect 235169 68147 235203 68175
rect 235231 68147 250377 68175
rect 250405 68147 250439 68175
rect 250467 68147 250501 68175
rect 250529 68147 250563 68175
rect 250591 68147 265737 68175
rect 265765 68147 265799 68175
rect 265827 68147 265861 68175
rect 265889 68147 265923 68175
rect 265951 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect -958 68113 298990 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 173577 68113
rect 173605 68085 173639 68113
rect 173667 68085 173701 68113
rect 173729 68085 173763 68113
rect 173791 68085 188937 68113
rect 188965 68085 188999 68113
rect 189027 68085 189061 68113
rect 189089 68085 189123 68113
rect 189151 68085 204297 68113
rect 204325 68085 204359 68113
rect 204387 68085 204421 68113
rect 204449 68085 204483 68113
rect 204511 68085 219657 68113
rect 219685 68085 219719 68113
rect 219747 68085 219781 68113
rect 219809 68085 219843 68113
rect 219871 68085 235017 68113
rect 235045 68085 235079 68113
rect 235107 68085 235141 68113
rect 235169 68085 235203 68113
rect 235231 68085 250377 68113
rect 250405 68085 250439 68113
rect 250467 68085 250501 68113
rect 250529 68085 250563 68113
rect 250591 68085 265737 68113
rect 265765 68085 265799 68113
rect 265827 68085 265861 68113
rect 265889 68085 265923 68113
rect 265951 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect -958 68051 298990 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 173577 68051
rect 173605 68023 173639 68051
rect 173667 68023 173701 68051
rect 173729 68023 173763 68051
rect 173791 68023 188937 68051
rect 188965 68023 188999 68051
rect 189027 68023 189061 68051
rect 189089 68023 189123 68051
rect 189151 68023 204297 68051
rect 204325 68023 204359 68051
rect 204387 68023 204421 68051
rect 204449 68023 204483 68051
rect 204511 68023 219657 68051
rect 219685 68023 219719 68051
rect 219747 68023 219781 68051
rect 219809 68023 219843 68051
rect 219871 68023 235017 68051
rect 235045 68023 235079 68051
rect 235107 68023 235141 68051
rect 235169 68023 235203 68051
rect 235231 68023 250377 68051
rect 250405 68023 250439 68051
rect 250467 68023 250501 68051
rect 250529 68023 250563 68051
rect 250591 68023 265737 68051
rect 265765 68023 265799 68051
rect 265827 68023 265861 68051
rect 265889 68023 265923 68051
rect 265951 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect -958 67989 298990 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 173577 67989
rect 173605 67961 173639 67989
rect 173667 67961 173701 67989
rect 173729 67961 173763 67989
rect 173791 67961 188937 67989
rect 188965 67961 188999 67989
rect 189027 67961 189061 67989
rect 189089 67961 189123 67989
rect 189151 67961 204297 67989
rect 204325 67961 204359 67989
rect 204387 67961 204421 67989
rect 204449 67961 204483 67989
rect 204511 67961 219657 67989
rect 219685 67961 219719 67989
rect 219747 67961 219781 67989
rect 219809 67961 219843 67989
rect 219871 67961 235017 67989
rect 235045 67961 235079 67989
rect 235107 67961 235141 67989
rect 235169 67961 235203 67989
rect 235231 67961 250377 67989
rect 250405 67961 250439 67989
rect 250467 67961 250501 67989
rect 250529 67961 250563 67989
rect 250591 67961 265737 67989
rect 265765 67961 265799 67989
rect 265827 67961 265861 67989
rect 265889 67961 265923 67989
rect 265951 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect -958 67913 298990 67961
rect -958 65175 298990 65223
rect -958 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 171717 65175
rect 171745 65147 171779 65175
rect 171807 65147 171841 65175
rect 171869 65147 171903 65175
rect 171931 65147 187077 65175
rect 187105 65147 187139 65175
rect 187167 65147 187201 65175
rect 187229 65147 187263 65175
rect 187291 65147 202437 65175
rect 202465 65147 202499 65175
rect 202527 65147 202561 65175
rect 202589 65147 202623 65175
rect 202651 65147 217797 65175
rect 217825 65147 217859 65175
rect 217887 65147 217921 65175
rect 217949 65147 217983 65175
rect 218011 65147 233157 65175
rect 233185 65147 233219 65175
rect 233247 65147 233281 65175
rect 233309 65147 233343 65175
rect 233371 65147 248517 65175
rect 248545 65147 248579 65175
rect 248607 65147 248641 65175
rect 248669 65147 248703 65175
rect 248731 65147 263877 65175
rect 263905 65147 263939 65175
rect 263967 65147 264001 65175
rect 264029 65147 264063 65175
rect 264091 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298990 65175
rect -958 65113 298990 65147
rect -958 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 171717 65113
rect 171745 65085 171779 65113
rect 171807 65085 171841 65113
rect 171869 65085 171903 65113
rect 171931 65085 187077 65113
rect 187105 65085 187139 65113
rect 187167 65085 187201 65113
rect 187229 65085 187263 65113
rect 187291 65085 202437 65113
rect 202465 65085 202499 65113
rect 202527 65085 202561 65113
rect 202589 65085 202623 65113
rect 202651 65085 217797 65113
rect 217825 65085 217859 65113
rect 217887 65085 217921 65113
rect 217949 65085 217983 65113
rect 218011 65085 233157 65113
rect 233185 65085 233219 65113
rect 233247 65085 233281 65113
rect 233309 65085 233343 65113
rect 233371 65085 248517 65113
rect 248545 65085 248579 65113
rect 248607 65085 248641 65113
rect 248669 65085 248703 65113
rect 248731 65085 263877 65113
rect 263905 65085 263939 65113
rect 263967 65085 264001 65113
rect 264029 65085 264063 65113
rect 264091 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298990 65113
rect -958 65051 298990 65085
rect -958 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 171717 65051
rect 171745 65023 171779 65051
rect 171807 65023 171841 65051
rect 171869 65023 171903 65051
rect 171931 65023 187077 65051
rect 187105 65023 187139 65051
rect 187167 65023 187201 65051
rect 187229 65023 187263 65051
rect 187291 65023 202437 65051
rect 202465 65023 202499 65051
rect 202527 65023 202561 65051
rect 202589 65023 202623 65051
rect 202651 65023 217797 65051
rect 217825 65023 217859 65051
rect 217887 65023 217921 65051
rect 217949 65023 217983 65051
rect 218011 65023 233157 65051
rect 233185 65023 233219 65051
rect 233247 65023 233281 65051
rect 233309 65023 233343 65051
rect 233371 65023 248517 65051
rect 248545 65023 248579 65051
rect 248607 65023 248641 65051
rect 248669 65023 248703 65051
rect 248731 65023 263877 65051
rect 263905 65023 263939 65051
rect 263967 65023 264001 65051
rect 264029 65023 264063 65051
rect 264091 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298990 65051
rect -958 64989 298990 65023
rect -958 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 171717 64989
rect 171745 64961 171779 64989
rect 171807 64961 171841 64989
rect 171869 64961 171903 64989
rect 171931 64961 187077 64989
rect 187105 64961 187139 64989
rect 187167 64961 187201 64989
rect 187229 64961 187263 64989
rect 187291 64961 202437 64989
rect 202465 64961 202499 64989
rect 202527 64961 202561 64989
rect 202589 64961 202623 64989
rect 202651 64961 217797 64989
rect 217825 64961 217859 64989
rect 217887 64961 217921 64989
rect 217949 64961 217983 64989
rect 218011 64961 233157 64989
rect 233185 64961 233219 64989
rect 233247 64961 233281 64989
rect 233309 64961 233343 64989
rect 233371 64961 248517 64989
rect 248545 64961 248579 64989
rect 248607 64961 248641 64989
rect 248669 64961 248703 64989
rect 248731 64961 263877 64989
rect 263905 64961 263939 64989
rect 263967 64961 264001 64989
rect 264029 64961 264063 64989
rect 264091 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298990 64989
rect -958 64913 298990 64961
rect -958 59175 298990 59223
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 173577 59175
rect 173605 59147 173639 59175
rect 173667 59147 173701 59175
rect 173729 59147 173763 59175
rect 173791 59147 188937 59175
rect 188965 59147 188999 59175
rect 189027 59147 189061 59175
rect 189089 59147 189123 59175
rect 189151 59147 204297 59175
rect 204325 59147 204359 59175
rect 204387 59147 204421 59175
rect 204449 59147 204483 59175
rect 204511 59147 219657 59175
rect 219685 59147 219719 59175
rect 219747 59147 219781 59175
rect 219809 59147 219843 59175
rect 219871 59147 235017 59175
rect 235045 59147 235079 59175
rect 235107 59147 235141 59175
rect 235169 59147 235203 59175
rect 235231 59147 250377 59175
rect 250405 59147 250439 59175
rect 250467 59147 250501 59175
rect 250529 59147 250563 59175
rect 250591 59147 265737 59175
rect 265765 59147 265799 59175
rect 265827 59147 265861 59175
rect 265889 59147 265923 59175
rect 265951 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect -958 59113 298990 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 173577 59113
rect 173605 59085 173639 59113
rect 173667 59085 173701 59113
rect 173729 59085 173763 59113
rect 173791 59085 188937 59113
rect 188965 59085 188999 59113
rect 189027 59085 189061 59113
rect 189089 59085 189123 59113
rect 189151 59085 204297 59113
rect 204325 59085 204359 59113
rect 204387 59085 204421 59113
rect 204449 59085 204483 59113
rect 204511 59085 219657 59113
rect 219685 59085 219719 59113
rect 219747 59085 219781 59113
rect 219809 59085 219843 59113
rect 219871 59085 235017 59113
rect 235045 59085 235079 59113
rect 235107 59085 235141 59113
rect 235169 59085 235203 59113
rect 235231 59085 250377 59113
rect 250405 59085 250439 59113
rect 250467 59085 250501 59113
rect 250529 59085 250563 59113
rect 250591 59085 265737 59113
rect 265765 59085 265799 59113
rect 265827 59085 265861 59113
rect 265889 59085 265923 59113
rect 265951 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect -958 59051 298990 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 173577 59051
rect 173605 59023 173639 59051
rect 173667 59023 173701 59051
rect 173729 59023 173763 59051
rect 173791 59023 188937 59051
rect 188965 59023 188999 59051
rect 189027 59023 189061 59051
rect 189089 59023 189123 59051
rect 189151 59023 204297 59051
rect 204325 59023 204359 59051
rect 204387 59023 204421 59051
rect 204449 59023 204483 59051
rect 204511 59023 219657 59051
rect 219685 59023 219719 59051
rect 219747 59023 219781 59051
rect 219809 59023 219843 59051
rect 219871 59023 235017 59051
rect 235045 59023 235079 59051
rect 235107 59023 235141 59051
rect 235169 59023 235203 59051
rect 235231 59023 250377 59051
rect 250405 59023 250439 59051
rect 250467 59023 250501 59051
rect 250529 59023 250563 59051
rect 250591 59023 265737 59051
rect 265765 59023 265799 59051
rect 265827 59023 265861 59051
rect 265889 59023 265923 59051
rect 265951 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect -958 58989 298990 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 173577 58989
rect 173605 58961 173639 58989
rect 173667 58961 173701 58989
rect 173729 58961 173763 58989
rect 173791 58961 188937 58989
rect 188965 58961 188999 58989
rect 189027 58961 189061 58989
rect 189089 58961 189123 58989
rect 189151 58961 204297 58989
rect 204325 58961 204359 58989
rect 204387 58961 204421 58989
rect 204449 58961 204483 58989
rect 204511 58961 219657 58989
rect 219685 58961 219719 58989
rect 219747 58961 219781 58989
rect 219809 58961 219843 58989
rect 219871 58961 235017 58989
rect 235045 58961 235079 58989
rect 235107 58961 235141 58989
rect 235169 58961 235203 58989
rect 235231 58961 250377 58989
rect 250405 58961 250439 58989
rect 250467 58961 250501 58989
rect 250529 58961 250563 58989
rect 250591 58961 265737 58989
rect 265765 58961 265799 58989
rect 265827 58961 265861 58989
rect 265889 58961 265923 58989
rect 265951 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect -958 58913 298990 58961
rect -958 56175 298990 56223
rect -958 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 171717 56175
rect 171745 56147 171779 56175
rect 171807 56147 171841 56175
rect 171869 56147 171903 56175
rect 171931 56147 187077 56175
rect 187105 56147 187139 56175
rect 187167 56147 187201 56175
rect 187229 56147 187263 56175
rect 187291 56147 202437 56175
rect 202465 56147 202499 56175
rect 202527 56147 202561 56175
rect 202589 56147 202623 56175
rect 202651 56147 217797 56175
rect 217825 56147 217859 56175
rect 217887 56147 217921 56175
rect 217949 56147 217983 56175
rect 218011 56147 233157 56175
rect 233185 56147 233219 56175
rect 233247 56147 233281 56175
rect 233309 56147 233343 56175
rect 233371 56147 248517 56175
rect 248545 56147 248579 56175
rect 248607 56147 248641 56175
rect 248669 56147 248703 56175
rect 248731 56147 263877 56175
rect 263905 56147 263939 56175
rect 263967 56147 264001 56175
rect 264029 56147 264063 56175
rect 264091 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298990 56175
rect -958 56113 298990 56147
rect -958 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 171717 56113
rect 171745 56085 171779 56113
rect 171807 56085 171841 56113
rect 171869 56085 171903 56113
rect 171931 56085 187077 56113
rect 187105 56085 187139 56113
rect 187167 56085 187201 56113
rect 187229 56085 187263 56113
rect 187291 56085 202437 56113
rect 202465 56085 202499 56113
rect 202527 56085 202561 56113
rect 202589 56085 202623 56113
rect 202651 56085 217797 56113
rect 217825 56085 217859 56113
rect 217887 56085 217921 56113
rect 217949 56085 217983 56113
rect 218011 56085 233157 56113
rect 233185 56085 233219 56113
rect 233247 56085 233281 56113
rect 233309 56085 233343 56113
rect 233371 56085 248517 56113
rect 248545 56085 248579 56113
rect 248607 56085 248641 56113
rect 248669 56085 248703 56113
rect 248731 56085 263877 56113
rect 263905 56085 263939 56113
rect 263967 56085 264001 56113
rect 264029 56085 264063 56113
rect 264091 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298990 56113
rect -958 56051 298990 56085
rect -958 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 171717 56051
rect 171745 56023 171779 56051
rect 171807 56023 171841 56051
rect 171869 56023 171903 56051
rect 171931 56023 187077 56051
rect 187105 56023 187139 56051
rect 187167 56023 187201 56051
rect 187229 56023 187263 56051
rect 187291 56023 202437 56051
rect 202465 56023 202499 56051
rect 202527 56023 202561 56051
rect 202589 56023 202623 56051
rect 202651 56023 217797 56051
rect 217825 56023 217859 56051
rect 217887 56023 217921 56051
rect 217949 56023 217983 56051
rect 218011 56023 233157 56051
rect 233185 56023 233219 56051
rect 233247 56023 233281 56051
rect 233309 56023 233343 56051
rect 233371 56023 248517 56051
rect 248545 56023 248579 56051
rect 248607 56023 248641 56051
rect 248669 56023 248703 56051
rect 248731 56023 263877 56051
rect 263905 56023 263939 56051
rect 263967 56023 264001 56051
rect 264029 56023 264063 56051
rect 264091 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298990 56051
rect -958 55989 298990 56023
rect -958 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 171717 55989
rect 171745 55961 171779 55989
rect 171807 55961 171841 55989
rect 171869 55961 171903 55989
rect 171931 55961 187077 55989
rect 187105 55961 187139 55989
rect 187167 55961 187201 55989
rect 187229 55961 187263 55989
rect 187291 55961 202437 55989
rect 202465 55961 202499 55989
rect 202527 55961 202561 55989
rect 202589 55961 202623 55989
rect 202651 55961 217797 55989
rect 217825 55961 217859 55989
rect 217887 55961 217921 55989
rect 217949 55961 217983 55989
rect 218011 55961 233157 55989
rect 233185 55961 233219 55989
rect 233247 55961 233281 55989
rect 233309 55961 233343 55989
rect 233371 55961 248517 55989
rect 248545 55961 248579 55989
rect 248607 55961 248641 55989
rect 248669 55961 248703 55989
rect 248731 55961 263877 55989
rect 263905 55961 263939 55989
rect 263967 55961 264001 55989
rect 264029 55961 264063 55989
rect 264091 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298990 55989
rect -958 55913 298990 55961
rect -958 50175 298990 50223
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 173577 50175
rect 173605 50147 173639 50175
rect 173667 50147 173701 50175
rect 173729 50147 173763 50175
rect 173791 50147 188937 50175
rect 188965 50147 188999 50175
rect 189027 50147 189061 50175
rect 189089 50147 189123 50175
rect 189151 50147 204297 50175
rect 204325 50147 204359 50175
rect 204387 50147 204421 50175
rect 204449 50147 204483 50175
rect 204511 50147 219657 50175
rect 219685 50147 219719 50175
rect 219747 50147 219781 50175
rect 219809 50147 219843 50175
rect 219871 50147 235017 50175
rect 235045 50147 235079 50175
rect 235107 50147 235141 50175
rect 235169 50147 235203 50175
rect 235231 50147 250377 50175
rect 250405 50147 250439 50175
rect 250467 50147 250501 50175
rect 250529 50147 250563 50175
rect 250591 50147 265737 50175
rect 265765 50147 265799 50175
rect 265827 50147 265861 50175
rect 265889 50147 265923 50175
rect 265951 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect -958 50113 298990 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 173577 50113
rect 173605 50085 173639 50113
rect 173667 50085 173701 50113
rect 173729 50085 173763 50113
rect 173791 50085 188937 50113
rect 188965 50085 188999 50113
rect 189027 50085 189061 50113
rect 189089 50085 189123 50113
rect 189151 50085 204297 50113
rect 204325 50085 204359 50113
rect 204387 50085 204421 50113
rect 204449 50085 204483 50113
rect 204511 50085 219657 50113
rect 219685 50085 219719 50113
rect 219747 50085 219781 50113
rect 219809 50085 219843 50113
rect 219871 50085 235017 50113
rect 235045 50085 235079 50113
rect 235107 50085 235141 50113
rect 235169 50085 235203 50113
rect 235231 50085 250377 50113
rect 250405 50085 250439 50113
rect 250467 50085 250501 50113
rect 250529 50085 250563 50113
rect 250591 50085 265737 50113
rect 265765 50085 265799 50113
rect 265827 50085 265861 50113
rect 265889 50085 265923 50113
rect 265951 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect -958 50051 298990 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 173577 50051
rect 173605 50023 173639 50051
rect 173667 50023 173701 50051
rect 173729 50023 173763 50051
rect 173791 50023 188937 50051
rect 188965 50023 188999 50051
rect 189027 50023 189061 50051
rect 189089 50023 189123 50051
rect 189151 50023 204297 50051
rect 204325 50023 204359 50051
rect 204387 50023 204421 50051
rect 204449 50023 204483 50051
rect 204511 50023 219657 50051
rect 219685 50023 219719 50051
rect 219747 50023 219781 50051
rect 219809 50023 219843 50051
rect 219871 50023 235017 50051
rect 235045 50023 235079 50051
rect 235107 50023 235141 50051
rect 235169 50023 235203 50051
rect 235231 50023 250377 50051
rect 250405 50023 250439 50051
rect 250467 50023 250501 50051
rect 250529 50023 250563 50051
rect 250591 50023 265737 50051
rect 265765 50023 265799 50051
rect 265827 50023 265861 50051
rect 265889 50023 265923 50051
rect 265951 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect -958 49989 298990 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 173577 49989
rect 173605 49961 173639 49989
rect 173667 49961 173701 49989
rect 173729 49961 173763 49989
rect 173791 49961 188937 49989
rect 188965 49961 188999 49989
rect 189027 49961 189061 49989
rect 189089 49961 189123 49989
rect 189151 49961 204297 49989
rect 204325 49961 204359 49989
rect 204387 49961 204421 49989
rect 204449 49961 204483 49989
rect 204511 49961 219657 49989
rect 219685 49961 219719 49989
rect 219747 49961 219781 49989
rect 219809 49961 219843 49989
rect 219871 49961 235017 49989
rect 235045 49961 235079 49989
rect 235107 49961 235141 49989
rect 235169 49961 235203 49989
rect 235231 49961 250377 49989
rect 250405 49961 250439 49989
rect 250467 49961 250501 49989
rect 250529 49961 250563 49989
rect 250591 49961 265737 49989
rect 265765 49961 265799 49989
rect 265827 49961 265861 49989
rect 265889 49961 265923 49989
rect 265951 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect -958 49913 298990 49961
rect -958 47175 298990 47223
rect -958 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 171717 47175
rect 171745 47147 171779 47175
rect 171807 47147 171841 47175
rect 171869 47147 171903 47175
rect 171931 47147 187077 47175
rect 187105 47147 187139 47175
rect 187167 47147 187201 47175
rect 187229 47147 187263 47175
rect 187291 47147 202437 47175
rect 202465 47147 202499 47175
rect 202527 47147 202561 47175
rect 202589 47147 202623 47175
rect 202651 47147 217797 47175
rect 217825 47147 217859 47175
rect 217887 47147 217921 47175
rect 217949 47147 217983 47175
rect 218011 47147 233157 47175
rect 233185 47147 233219 47175
rect 233247 47147 233281 47175
rect 233309 47147 233343 47175
rect 233371 47147 248517 47175
rect 248545 47147 248579 47175
rect 248607 47147 248641 47175
rect 248669 47147 248703 47175
rect 248731 47147 263877 47175
rect 263905 47147 263939 47175
rect 263967 47147 264001 47175
rect 264029 47147 264063 47175
rect 264091 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298990 47175
rect -958 47113 298990 47147
rect -958 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 171717 47113
rect 171745 47085 171779 47113
rect 171807 47085 171841 47113
rect 171869 47085 171903 47113
rect 171931 47085 187077 47113
rect 187105 47085 187139 47113
rect 187167 47085 187201 47113
rect 187229 47085 187263 47113
rect 187291 47085 202437 47113
rect 202465 47085 202499 47113
rect 202527 47085 202561 47113
rect 202589 47085 202623 47113
rect 202651 47085 217797 47113
rect 217825 47085 217859 47113
rect 217887 47085 217921 47113
rect 217949 47085 217983 47113
rect 218011 47085 233157 47113
rect 233185 47085 233219 47113
rect 233247 47085 233281 47113
rect 233309 47085 233343 47113
rect 233371 47085 248517 47113
rect 248545 47085 248579 47113
rect 248607 47085 248641 47113
rect 248669 47085 248703 47113
rect 248731 47085 263877 47113
rect 263905 47085 263939 47113
rect 263967 47085 264001 47113
rect 264029 47085 264063 47113
rect 264091 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298990 47113
rect -958 47051 298990 47085
rect -958 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 171717 47051
rect 171745 47023 171779 47051
rect 171807 47023 171841 47051
rect 171869 47023 171903 47051
rect 171931 47023 187077 47051
rect 187105 47023 187139 47051
rect 187167 47023 187201 47051
rect 187229 47023 187263 47051
rect 187291 47023 202437 47051
rect 202465 47023 202499 47051
rect 202527 47023 202561 47051
rect 202589 47023 202623 47051
rect 202651 47023 217797 47051
rect 217825 47023 217859 47051
rect 217887 47023 217921 47051
rect 217949 47023 217983 47051
rect 218011 47023 233157 47051
rect 233185 47023 233219 47051
rect 233247 47023 233281 47051
rect 233309 47023 233343 47051
rect 233371 47023 248517 47051
rect 248545 47023 248579 47051
rect 248607 47023 248641 47051
rect 248669 47023 248703 47051
rect 248731 47023 263877 47051
rect 263905 47023 263939 47051
rect 263967 47023 264001 47051
rect 264029 47023 264063 47051
rect 264091 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298990 47051
rect -958 46989 298990 47023
rect -958 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 171717 46989
rect 171745 46961 171779 46989
rect 171807 46961 171841 46989
rect 171869 46961 171903 46989
rect 171931 46961 187077 46989
rect 187105 46961 187139 46989
rect 187167 46961 187201 46989
rect 187229 46961 187263 46989
rect 187291 46961 202437 46989
rect 202465 46961 202499 46989
rect 202527 46961 202561 46989
rect 202589 46961 202623 46989
rect 202651 46961 217797 46989
rect 217825 46961 217859 46989
rect 217887 46961 217921 46989
rect 217949 46961 217983 46989
rect 218011 46961 233157 46989
rect 233185 46961 233219 46989
rect 233247 46961 233281 46989
rect 233309 46961 233343 46989
rect 233371 46961 248517 46989
rect 248545 46961 248579 46989
rect 248607 46961 248641 46989
rect 248669 46961 248703 46989
rect 248731 46961 263877 46989
rect 263905 46961 263939 46989
rect 263967 46961 264001 46989
rect 264029 46961 264063 46989
rect 264091 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298990 46989
rect -958 46913 298990 46961
rect -958 41175 298990 41223
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 173577 41175
rect 173605 41147 173639 41175
rect 173667 41147 173701 41175
rect 173729 41147 173763 41175
rect 173791 41147 188937 41175
rect 188965 41147 188999 41175
rect 189027 41147 189061 41175
rect 189089 41147 189123 41175
rect 189151 41147 204297 41175
rect 204325 41147 204359 41175
rect 204387 41147 204421 41175
rect 204449 41147 204483 41175
rect 204511 41147 219657 41175
rect 219685 41147 219719 41175
rect 219747 41147 219781 41175
rect 219809 41147 219843 41175
rect 219871 41147 235017 41175
rect 235045 41147 235079 41175
rect 235107 41147 235141 41175
rect 235169 41147 235203 41175
rect 235231 41147 250377 41175
rect 250405 41147 250439 41175
rect 250467 41147 250501 41175
rect 250529 41147 250563 41175
rect 250591 41147 265737 41175
rect 265765 41147 265799 41175
rect 265827 41147 265861 41175
rect 265889 41147 265923 41175
rect 265951 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect -958 41113 298990 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 173577 41113
rect 173605 41085 173639 41113
rect 173667 41085 173701 41113
rect 173729 41085 173763 41113
rect 173791 41085 188937 41113
rect 188965 41085 188999 41113
rect 189027 41085 189061 41113
rect 189089 41085 189123 41113
rect 189151 41085 204297 41113
rect 204325 41085 204359 41113
rect 204387 41085 204421 41113
rect 204449 41085 204483 41113
rect 204511 41085 219657 41113
rect 219685 41085 219719 41113
rect 219747 41085 219781 41113
rect 219809 41085 219843 41113
rect 219871 41085 235017 41113
rect 235045 41085 235079 41113
rect 235107 41085 235141 41113
rect 235169 41085 235203 41113
rect 235231 41085 250377 41113
rect 250405 41085 250439 41113
rect 250467 41085 250501 41113
rect 250529 41085 250563 41113
rect 250591 41085 265737 41113
rect 265765 41085 265799 41113
rect 265827 41085 265861 41113
rect 265889 41085 265923 41113
rect 265951 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect -958 41051 298990 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 173577 41051
rect 173605 41023 173639 41051
rect 173667 41023 173701 41051
rect 173729 41023 173763 41051
rect 173791 41023 188937 41051
rect 188965 41023 188999 41051
rect 189027 41023 189061 41051
rect 189089 41023 189123 41051
rect 189151 41023 204297 41051
rect 204325 41023 204359 41051
rect 204387 41023 204421 41051
rect 204449 41023 204483 41051
rect 204511 41023 219657 41051
rect 219685 41023 219719 41051
rect 219747 41023 219781 41051
rect 219809 41023 219843 41051
rect 219871 41023 235017 41051
rect 235045 41023 235079 41051
rect 235107 41023 235141 41051
rect 235169 41023 235203 41051
rect 235231 41023 250377 41051
rect 250405 41023 250439 41051
rect 250467 41023 250501 41051
rect 250529 41023 250563 41051
rect 250591 41023 265737 41051
rect 265765 41023 265799 41051
rect 265827 41023 265861 41051
rect 265889 41023 265923 41051
rect 265951 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect -958 40989 298990 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 173577 40989
rect 173605 40961 173639 40989
rect 173667 40961 173701 40989
rect 173729 40961 173763 40989
rect 173791 40961 188937 40989
rect 188965 40961 188999 40989
rect 189027 40961 189061 40989
rect 189089 40961 189123 40989
rect 189151 40961 204297 40989
rect 204325 40961 204359 40989
rect 204387 40961 204421 40989
rect 204449 40961 204483 40989
rect 204511 40961 219657 40989
rect 219685 40961 219719 40989
rect 219747 40961 219781 40989
rect 219809 40961 219843 40989
rect 219871 40961 235017 40989
rect 235045 40961 235079 40989
rect 235107 40961 235141 40989
rect 235169 40961 235203 40989
rect 235231 40961 250377 40989
rect 250405 40961 250439 40989
rect 250467 40961 250501 40989
rect 250529 40961 250563 40989
rect 250591 40961 265737 40989
rect 265765 40961 265799 40989
rect 265827 40961 265861 40989
rect 265889 40961 265923 40989
rect 265951 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect -958 40913 298990 40961
rect -958 38175 298990 38223
rect -958 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 171717 38175
rect 171745 38147 171779 38175
rect 171807 38147 171841 38175
rect 171869 38147 171903 38175
rect 171931 38147 187077 38175
rect 187105 38147 187139 38175
rect 187167 38147 187201 38175
rect 187229 38147 187263 38175
rect 187291 38147 202437 38175
rect 202465 38147 202499 38175
rect 202527 38147 202561 38175
rect 202589 38147 202623 38175
rect 202651 38147 217797 38175
rect 217825 38147 217859 38175
rect 217887 38147 217921 38175
rect 217949 38147 217983 38175
rect 218011 38147 233157 38175
rect 233185 38147 233219 38175
rect 233247 38147 233281 38175
rect 233309 38147 233343 38175
rect 233371 38147 248517 38175
rect 248545 38147 248579 38175
rect 248607 38147 248641 38175
rect 248669 38147 248703 38175
rect 248731 38147 263877 38175
rect 263905 38147 263939 38175
rect 263967 38147 264001 38175
rect 264029 38147 264063 38175
rect 264091 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298990 38175
rect -958 38113 298990 38147
rect -958 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 171717 38113
rect 171745 38085 171779 38113
rect 171807 38085 171841 38113
rect 171869 38085 171903 38113
rect 171931 38085 187077 38113
rect 187105 38085 187139 38113
rect 187167 38085 187201 38113
rect 187229 38085 187263 38113
rect 187291 38085 202437 38113
rect 202465 38085 202499 38113
rect 202527 38085 202561 38113
rect 202589 38085 202623 38113
rect 202651 38085 217797 38113
rect 217825 38085 217859 38113
rect 217887 38085 217921 38113
rect 217949 38085 217983 38113
rect 218011 38085 233157 38113
rect 233185 38085 233219 38113
rect 233247 38085 233281 38113
rect 233309 38085 233343 38113
rect 233371 38085 248517 38113
rect 248545 38085 248579 38113
rect 248607 38085 248641 38113
rect 248669 38085 248703 38113
rect 248731 38085 263877 38113
rect 263905 38085 263939 38113
rect 263967 38085 264001 38113
rect 264029 38085 264063 38113
rect 264091 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298990 38113
rect -958 38051 298990 38085
rect -958 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 171717 38051
rect 171745 38023 171779 38051
rect 171807 38023 171841 38051
rect 171869 38023 171903 38051
rect 171931 38023 187077 38051
rect 187105 38023 187139 38051
rect 187167 38023 187201 38051
rect 187229 38023 187263 38051
rect 187291 38023 202437 38051
rect 202465 38023 202499 38051
rect 202527 38023 202561 38051
rect 202589 38023 202623 38051
rect 202651 38023 217797 38051
rect 217825 38023 217859 38051
rect 217887 38023 217921 38051
rect 217949 38023 217983 38051
rect 218011 38023 233157 38051
rect 233185 38023 233219 38051
rect 233247 38023 233281 38051
rect 233309 38023 233343 38051
rect 233371 38023 248517 38051
rect 248545 38023 248579 38051
rect 248607 38023 248641 38051
rect 248669 38023 248703 38051
rect 248731 38023 263877 38051
rect 263905 38023 263939 38051
rect 263967 38023 264001 38051
rect 264029 38023 264063 38051
rect 264091 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298990 38051
rect -958 37989 298990 38023
rect -958 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 171717 37989
rect 171745 37961 171779 37989
rect 171807 37961 171841 37989
rect 171869 37961 171903 37989
rect 171931 37961 187077 37989
rect 187105 37961 187139 37989
rect 187167 37961 187201 37989
rect 187229 37961 187263 37989
rect 187291 37961 202437 37989
rect 202465 37961 202499 37989
rect 202527 37961 202561 37989
rect 202589 37961 202623 37989
rect 202651 37961 217797 37989
rect 217825 37961 217859 37989
rect 217887 37961 217921 37989
rect 217949 37961 217983 37989
rect 218011 37961 233157 37989
rect 233185 37961 233219 37989
rect 233247 37961 233281 37989
rect 233309 37961 233343 37989
rect 233371 37961 248517 37989
rect 248545 37961 248579 37989
rect 248607 37961 248641 37989
rect 248669 37961 248703 37989
rect 248731 37961 263877 37989
rect 263905 37961 263939 37989
rect 263967 37961 264001 37989
rect 264029 37961 264063 37989
rect 264091 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298990 37989
rect -958 37913 298990 37961
rect -958 32175 298990 32223
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 173577 32175
rect 173605 32147 173639 32175
rect 173667 32147 173701 32175
rect 173729 32147 173763 32175
rect 173791 32147 188937 32175
rect 188965 32147 188999 32175
rect 189027 32147 189061 32175
rect 189089 32147 189123 32175
rect 189151 32147 204297 32175
rect 204325 32147 204359 32175
rect 204387 32147 204421 32175
rect 204449 32147 204483 32175
rect 204511 32147 219657 32175
rect 219685 32147 219719 32175
rect 219747 32147 219781 32175
rect 219809 32147 219843 32175
rect 219871 32147 235017 32175
rect 235045 32147 235079 32175
rect 235107 32147 235141 32175
rect 235169 32147 235203 32175
rect 235231 32147 250377 32175
rect 250405 32147 250439 32175
rect 250467 32147 250501 32175
rect 250529 32147 250563 32175
rect 250591 32147 265737 32175
rect 265765 32147 265799 32175
rect 265827 32147 265861 32175
rect 265889 32147 265923 32175
rect 265951 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect -958 32113 298990 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 173577 32113
rect 173605 32085 173639 32113
rect 173667 32085 173701 32113
rect 173729 32085 173763 32113
rect 173791 32085 188937 32113
rect 188965 32085 188999 32113
rect 189027 32085 189061 32113
rect 189089 32085 189123 32113
rect 189151 32085 204297 32113
rect 204325 32085 204359 32113
rect 204387 32085 204421 32113
rect 204449 32085 204483 32113
rect 204511 32085 219657 32113
rect 219685 32085 219719 32113
rect 219747 32085 219781 32113
rect 219809 32085 219843 32113
rect 219871 32085 235017 32113
rect 235045 32085 235079 32113
rect 235107 32085 235141 32113
rect 235169 32085 235203 32113
rect 235231 32085 250377 32113
rect 250405 32085 250439 32113
rect 250467 32085 250501 32113
rect 250529 32085 250563 32113
rect 250591 32085 265737 32113
rect 265765 32085 265799 32113
rect 265827 32085 265861 32113
rect 265889 32085 265923 32113
rect 265951 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect -958 32051 298990 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 173577 32051
rect 173605 32023 173639 32051
rect 173667 32023 173701 32051
rect 173729 32023 173763 32051
rect 173791 32023 188937 32051
rect 188965 32023 188999 32051
rect 189027 32023 189061 32051
rect 189089 32023 189123 32051
rect 189151 32023 204297 32051
rect 204325 32023 204359 32051
rect 204387 32023 204421 32051
rect 204449 32023 204483 32051
rect 204511 32023 219657 32051
rect 219685 32023 219719 32051
rect 219747 32023 219781 32051
rect 219809 32023 219843 32051
rect 219871 32023 235017 32051
rect 235045 32023 235079 32051
rect 235107 32023 235141 32051
rect 235169 32023 235203 32051
rect 235231 32023 250377 32051
rect 250405 32023 250439 32051
rect 250467 32023 250501 32051
rect 250529 32023 250563 32051
rect 250591 32023 265737 32051
rect 265765 32023 265799 32051
rect 265827 32023 265861 32051
rect 265889 32023 265923 32051
rect 265951 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect -958 31989 298990 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 173577 31989
rect 173605 31961 173639 31989
rect 173667 31961 173701 31989
rect 173729 31961 173763 31989
rect 173791 31961 188937 31989
rect 188965 31961 188999 31989
rect 189027 31961 189061 31989
rect 189089 31961 189123 31989
rect 189151 31961 204297 31989
rect 204325 31961 204359 31989
rect 204387 31961 204421 31989
rect 204449 31961 204483 31989
rect 204511 31961 219657 31989
rect 219685 31961 219719 31989
rect 219747 31961 219781 31989
rect 219809 31961 219843 31989
rect 219871 31961 235017 31989
rect 235045 31961 235079 31989
rect 235107 31961 235141 31989
rect 235169 31961 235203 31989
rect 235231 31961 250377 31989
rect 250405 31961 250439 31989
rect 250467 31961 250501 31989
rect 250529 31961 250563 31989
rect 250591 31961 265737 31989
rect 265765 31961 265799 31989
rect 265827 31961 265861 31989
rect 265889 31961 265923 31989
rect 265951 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect -958 31913 298990 31961
rect -958 29175 298990 29223
rect -958 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 171717 29175
rect 171745 29147 171779 29175
rect 171807 29147 171841 29175
rect 171869 29147 171903 29175
rect 171931 29147 187077 29175
rect 187105 29147 187139 29175
rect 187167 29147 187201 29175
rect 187229 29147 187263 29175
rect 187291 29147 202437 29175
rect 202465 29147 202499 29175
rect 202527 29147 202561 29175
rect 202589 29147 202623 29175
rect 202651 29147 217797 29175
rect 217825 29147 217859 29175
rect 217887 29147 217921 29175
rect 217949 29147 217983 29175
rect 218011 29147 233157 29175
rect 233185 29147 233219 29175
rect 233247 29147 233281 29175
rect 233309 29147 233343 29175
rect 233371 29147 248517 29175
rect 248545 29147 248579 29175
rect 248607 29147 248641 29175
rect 248669 29147 248703 29175
rect 248731 29147 263877 29175
rect 263905 29147 263939 29175
rect 263967 29147 264001 29175
rect 264029 29147 264063 29175
rect 264091 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298990 29175
rect -958 29113 298990 29147
rect -958 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 171717 29113
rect 171745 29085 171779 29113
rect 171807 29085 171841 29113
rect 171869 29085 171903 29113
rect 171931 29085 187077 29113
rect 187105 29085 187139 29113
rect 187167 29085 187201 29113
rect 187229 29085 187263 29113
rect 187291 29085 202437 29113
rect 202465 29085 202499 29113
rect 202527 29085 202561 29113
rect 202589 29085 202623 29113
rect 202651 29085 217797 29113
rect 217825 29085 217859 29113
rect 217887 29085 217921 29113
rect 217949 29085 217983 29113
rect 218011 29085 233157 29113
rect 233185 29085 233219 29113
rect 233247 29085 233281 29113
rect 233309 29085 233343 29113
rect 233371 29085 248517 29113
rect 248545 29085 248579 29113
rect 248607 29085 248641 29113
rect 248669 29085 248703 29113
rect 248731 29085 263877 29113
rect 263905 29085 263939 29113
rect 263967 29085 264001 29113
rect 264029 29085 264063 29113
rect 264091 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298990 29113
rect -958 29051 298990 29085
rect -958 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 171717 29051
rect 171745 29023 171779 29051
rect 171807 29023 171841 29051
rect 171869 29023 171903 29051
rect 171931 29023 187077 29051
rect 187105 29023 187139 29051
rect 187167 29023 187201 29051
rect 187229 29023 187263 29051
rect 187291 29023 202437 29051
rect 202465 29023 202499 29051
rect 202527 29023 202561 29051
rect 202589 29023 202623 29051
rect 202651 29023 217797 29051
rect 217825 29023 217859 29051
rect 217887 29023 217921 29051
rect 217949 29023 217983 29051
rect 218011 29023 233157 29051
rect 233185 29023 233219 29051
rect 233247 29023 233281 29051
rect 233309 29023 233343 29051
rect 233371 29023 248517 29051
rect 248545 29023 248579 29051
rect 248607 29023 248641 29051
rect 248669 29023 248703 29051
rect 248731 29023 263877 29051
rect 263905 29023 263939 29051
rect 263967 29023 264001 29051
rect 264029 29023 264063 29051
rect 264091 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298990 29051
rect -958 28989 298990 29023
rect -958 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 171717 28989
rect 171745 28961 171779 28989
rect 171807 28961 171841 28989
rect 171869 28961 171903 28989
rect 171931 28961 187077 28989
rect 187105 28961 187139 28989
rect 187167 28961 187201 28989
rect 187229 28961 187263 28989
rect 187291 28961 202437 28989
rect 202465 28961 202499 28989
rect 202527 28961 202561 28989
rect 202589 28961 202623 28989
rect 202651 28961 217797 28989
rect 217825 28961 217859 28989
rect 217887 28961 217921 28989
rect 217949 28961 217983 28989
rect 218011 28961 233157 28989
rect 233185 28961 233219 28989
rect 233247 28961 233281 28989
rect 233309 28961 233343 28989
rect 233371 28961 248517 28989
rect 248545 28961 248579 28989
rect 248607 28961 248641 28989
rect 248669 28961 248703 28989
rect 248731 28961 263877 28989
rect 263905 28961 263939 28989
rect 263967 28961 264001 28989
rect 264029 28961 264063 28989
rect 264091 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298990 28989
rect -958 28913 298990 28961
rect -958 23175 298990 23223
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 173577 23175
rect 173605 23147 173639 23175
rect 173667 23147 173701 23175
rect 173729 23147 173763 23175
rect 173791 23147 188937 23175
rect 188965 23147 188999 23175
rect 189027 23147 189061 23175
rect 189089 23147 189123 23175
rect 189151 23147 204297 23175
rect 204325 23147 204359 23175
rect 204387 23147 204421 23175
rect 204449 23147 204483 23175
rect 204511 23147 219657 23175
rect 219685 23147 219719 23175
rect 219747 23147 219781 23175
rect 219809 23147 219843 23175
rect 219871 23147 235017 23175
rect 235045 23147 235079 23175
rect 235107 23147 235141 23175
rect 235169 23147 235203 23175
rect 235231 23147 250377 23175
rect 250405 23147 250439 23175
rect 250467 23147 250501 23175
rect 250529 23147 250563 23175
rect 250591 23147 265737 23175
rect 265765 23147 265799 23175
rect 265827 23147 265861 23175
rect 265889 23147 265923 23175
rect 265951 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect -958 23113 298990 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 173577 23113
rect 173605 23085 173639 23113
rect 173667 23085 173701 23113
rect 173729 23085 173763 23113
rect 173791 23085 188937 23113
rect 188965 23085 188999 23113
rect 189027 23085 189061 23113
rect 189089 23085 189123 23113
rect 189151 23085 204297 23113
rect 204325 23085 204359 23113
rect 204387 23085 204421 23113
rect 204449 23085 204483 23113
rect 204511 23085 219657 23113
rect 219685 23085 219719 23113
rect 219747 23085 219781 23113
rect 219809 23085 219843 23113
rect 219871 23085 235017 23113
rect 235045 23085 235079 23113
rect 235107 23085 235141 23113
rect 235169 23085 235203 23113
rect 235231 23085 250377 23113
rect 250405 23085 250439 23113
rect 250467 23085 250501 23113
rect 250529 23085 250563 23113
rect 250591 23085 265737 23113
rect 265765 23085 265799 23113
rect 265827 23085 265861 23113
rect 265889 23085 265923 23113
rect 265951 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect -958 23051 298990 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 173577 23051
rect 173605 23023 173639 23051
rect 173667 23023 173701 23051
rect 173729 23023 173763 23051
rect 173791 23023 188937 23051
rect 188965 23023 188999 23051
rect 189027 23023 189061 23051
rect 189089 23023 189123 23051
rect 189151 23023 204297 23051
rect 204325 23023 204359 23051
rect 204387 23023 204421 23051
rect 204449 23023 204483 23051
rect 204511 23023 219657 23051
rect 219685 23023 219719 23051
rect 219747 23023 219781 23051
rect 219809 23023 219843 23051
rect 219871 23023 235017 23051
rect 235045 23023 235079 23051
rect 235107 23023 235141 23051
rect 235169 23023 235203 23051
rect 235231 23023 250377 23051
rect 250405 23023 250439 23051
rect 250467 23023 250501 23051
rect 250529 23023 250563 23051
rect 250591 23023 265737 23051
rect 265765 23023 265799 23051
rect 265827 23023 265861 23051
rect 265889 23023 265923 23051
rect 265951 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect -958 22989 298990 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 173577 22989
rect 173605 22961 173639 22989
rect 173667 22961 173701 22989
rect 173729 22961 173763 22989
rect 173791 22961 188937 22989
rect 188965 22961 188999 22989
rect 189027 22961 189061 22989
rect 189089 22961 189123 22989
rect 189151 22961 204297 22989
rect 204325 22961 204359 22989
rect 204387 22961 204421 22989
rect 204449 22961 204483 22989
rect 204511 22961 219657 22989
rect 219685 22961 219719 22989
rect 219747 22961 219781 22989
rect 219809 22961 219843 22989
rect 219871 22961 235017 22989
rect 235045 22961 235079 22989
rect 235107 22961 235141 22989
rect 235169 22961 235203 22989
rect 235231 22961 250377 22989
rect 250405 22961 250439 22989
rect 250467 22961 250501 22989
rect 250529 22961 250563 22989
rect 250591 22961 265737 22989
rect 265765 22961 265799 22989
rect 265827 22961 265861 22989
rect 265889 22961 265923 22989
rect 265951 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect -958 22913 298990 22961
rect -958 20175 298990 20223
rect -958 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 171717 20175
rect 171745 20147 171779 20175
rect 171807 20147 171841 20175
rect 171869 20147 171903 20175
rect 171931 20147 187077 20175
rect 187105 20147 187139 20175
rect 187167 20147 187201 20175
rect 187229 20147 187263 20175
rect 187291 20147 202437 20175
rect 202465 20147 202499 20175
rect 202527 20147 202561 20175
rect 202589 20147 202623 20175
rect 202651 20147 217797 20175
rect 217825 20147 217859 20175
rect 217887 20147 217921 20175
rect 217949 20147 217983 20175
rect 218011 20147 233157 20175
rect 233185 20147 233219 20175
rect 233247 20147 233281 20175
rect 233309 20147 233343 20175
rect 233371 20147 248517 20175
rect 248545 20147 248579 20175
rect 248607 20147 248641 20175
rect 248669 20147 248703 20175
rect 248731 20147 263877 20175
rect 263905 20147 263939 20175
rect 263967 20147 264001 20175
rect 264029 20147 264063 20175
rect 264091 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298990 20175
rect -958 20113 298990 20147
rect -958 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 171717 20113
rect 171745 20085 171779 20113
rect 171807 20085 171841 20113
rect 171869 20085 171903 20113
rect 171931 20085 187077 20113
rect 187105 20085 187139 20113
rect 187167 20085 187201 20113
rect 187229 20085 187263 20113
rect 187291 20085 202437 20113
rect 202465 20085 202499 20113
rect 202527 20085 202561 20113
rect 202589 20085 202623 20113
rect 202651 20085 217797 20113
rect 217825 20085 217859 20113
rect 217887 20085 217921 20113
rect 217949 20085 217983 20113
rect 218011 20085 233157 20113
rect 233185 20085 233219 20113
rect 233247 20085 233281 20113
rect 233309 20085 233343 20113
rect 233371 20085 248517 20113
rect 248545 20085 248579 20113
rect 248607 20085 248641 20113
rect 248669 20085 248703 20113
rect 248731 20085 263877 20113
rect 263905 20085 263939 20113
rect 263967 20085 264001 20113
rect 264029 20085 264063 20113
rect 264091 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298990 20113
rect -958 20051 298990 20085
rect -958 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 171717 20051
rect 171745 20023 171779 20051
rect 171807 20023 171841 20051
rect 171869 20023 171903 20051
rect 171931 20023 187077 20051
rect 187105 20023 187139 20051
rect 187167 20023 187201 20051
rect 187229 20023 187263 20051
rect 187291 20023 202437 20051
rect 202465 20023 202499 20051
rect 202527 20023 202561 20051
rect 202589 20023 202623 20051
rect 202651 20023 217797 20051
rect 217825 20023 217859 20051
rect 217887 20023 217921 20051
rect 217949 20023 217983 20051
rect 218011 20023 233157 20051
rect 233185 20023 233219 20051
rect 233247 20023 233281 20051
rect 233309 20023 233343 20051
rect 233371 20023 248517 20051
rect 248545 20023 248579 20051
rect 248607 20023 248641 20051
rect 248669 20023 248703 20051
rect 248731 20023 263877 20051
rect 263905 20023 263939 20051
rect 263967 20023 264001 20051
rect 264029 20023 264063 20051
rect 264091 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298990 20051
rect -958 19989 298990 20023
rect -958 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 171717 19989
rect 171745 19961 171779 19989
rect 171807 19961 171841 19989
rect 171869 19961 171903 19989
rect 171931 19961 187077 19989
rect 187105 19961 187139 19989
rect 187167 19961 187201 19989
rect 187229 19961 187263 19989
rect 187291 19961 202437 19989
rect 202465 19961 202499 19989
rect 202527 19961 202561 19989
rect 202589 19961 202623 19989
rect 202651 19961 217797 19989
rect 217825 19961 217859 19989
rect 217887 19961 217921 19989
rect 217949 19961 217983 19989
rect 218011 19961 233157 19989
rect 233185 19961 233219 19989
rect 233247 19961 233281 19989
rect 233309 19961 233343 19989
rect 233371 19961 248517 19989
rect 248545 19961 248579 19989
rect 248607 19961 248641 19989
rect 248669 19961 248703 19989
rect 248731 19961 263877 19989
rect 263905 19961 263939 19989
rect 263967 19961 264001 19989
rect 264029 19961 264063 19989
rect 264091 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298990 19989
rect -958 19913 298990 19961
rect -958 14175 298990 14223
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 173577 14175
rect 173605 14147 173639 14175
rect 173667 14147 173701 14175
rect 173729 14147 173763 14175
rect 173791 14147 188937 14175
rect 188965 14147 188999 14175
rect 189027 14147 189061 14175
rect 189089 14147 189123 14175
rect 189151 14147 204297 14175
rect 204325 14147 204359 14175
rect 204387 14147 204421 14175
rect 204449 14147 204483 14175
rect 204511 14147 219657 14175
rect 219685 14147 219719 14175
rect 219747 14147 219781 14175
rect 219809 14147 219843 14175
rect 219871 14147 235017 14175
rect 235045 14147 235079 14175
rect 235107 14147 235141 14175
rect 235169 14147 235203 14175
rect 235231 14147 250377 14175
rect 250405 14147 250439 14175
rect 250467 14147 250501 14175
rect 250529 14147 250563 14175
rect 250591 14147 265737 14175
rect 265765 14147 265799 14175
rect 265827 14147 265861 14175
rect 265889 14147 265923 14175
rect 265951 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect -958 14113 298990 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 173577 14113
rect 173605 14085 173639 14113
rect 173667 14085 173701 14113
rect 173729 14085 173763 14113
rect 173791 14085 188937 14113
rect 188965 14085 188999 14113
rect 189027 14085 189061 14113
rect 189089 14085 189123 14113
rect 189151 14085 204297 14113
rect 204325 14085 204359 14113
rect 204387 14085 204421 14113
rect 204449 14085 204483 14113
rect 204511 14085 219657 14113
rect 219685 14085 219719 14113
rect 219747 14085 219781 14113
rect 219809 14085 219843 14113
rect 219871 14085 235017 14113
rect 235045 14085 235079 14113
rect 235107 14085 235141 14113
rect 235169 14085 235203 14113
rect 235231 14085 250377 14113
rect 250405 14085 250439 14113
rect 250467 14085 250501 14113
rect 250529 14085 250563 14113
rect 250591 14085 265737 14113
rect 265765 14085 265799 14113
rect 265827 14085 265861 14113
rect 265889 14085 265923 14113
rect 265951 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect -958 14051 298990 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 173577 14051
rect 173605 14023 173639 14051
rect 173667 14023 173701 14051
rect 173729 14023 173763 14051
rect 173791 14023 188937 14051
rect 188965 14023 188999 14051
rect 189027 14023 189061 14051
rect 189089 14023 189123 14051
rect 189151 14023 204297 14051
rect 204325 14023 204359 14051
rect 204387 14023 204421 14051
rect 204449 14023 204483 14051
rect 204511 14023 219657 14051
rect 219685 14023 219719 14051
rect 219747 14023 219781 14051
rect 219809 14023 219843 14051
rect 219871 14023 235017 14051
rect 235045 14023 235079 14051
rect 235107 14023 235141 14051
rect 235169 14023 235203 14051
rect 235231 14023 250377 14051
rect 250405 14023 250439 14051
rect 250467 14023 250501 14051
rect 250529 14023 250563 14051
rect 250591 14023 265737 14051
rect 265765 14023 265799 14051
rect 265827 14023 265861 14051
rect 265889 14023 265923 14051
rect 265951 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect -958 13989 298990 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 173577 13989
rect 173605 13961 173639 13989
rect 173667 13961 173701 13989
rect 173729 13961 173763 13989
rect 173791 13961 188937 13989
rect 188965 13961 188999 13989
rect 189027 13961 189061 13989
rect 189089 13961 189123 13989
rect 189151 13961 204297 13989
rect 204325 13961 204359 13989
rect 204387 13961 204421 13989
rect 204449 13961 204483 13989
rect 204511 13961 219657 13989
rect 219685 13961 219719 13989
rect 219747 13961 219781 13989
rect 219809 13961 219843 13989
rect 219871 13961 235017 13989
rect 235045 13961 235079 13989
rect 235107 13961 235141 13989
rect 235169 13961 235203 13989
rect 235231 13961 250377 13989
rect 250405 13961 250439 13989
rect 250467 13961 250501 13989
rect 250529 13961 250563 13989
rect 250591 13961 265737 13989
rect 265765 13961 265799 13989
rect 265827 13961 265861 13989
rect 265889 13961 265923 13989
rect 265951 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect -958 13913 298990 13961
rect -958 11175 298990 11223
rect -958 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 171717 11175
rect 171745 11147 171779 11175
rect 171807 11147 171841 11175
rect 171869 11147 171903 11175
rect 171931 11147 187077 11175
rect 187105 11147 187139 11175
rect 187167 11147 187201 11175
rect 187229 11147 187263 11175
rect 187291 11147 202437 11175
rect 202465 11147 202499 11175
rect 202527 11147 202561 11175
rect 202589 11147 202623 11175
rect 202651 11147 217797 11175
rect 217825 11147 217859 11175
rect 217887 11147 217921 11175
rect 217949 11147 217983 11175
rect 218011 11147 233157 11175
rect 233185 11147 233219 11175
rect 233247 11147 233281 11175
rect 233309 11147 233343 11175
rect 233371 11147 248517 11175
rect 248545 11147 248579 11175
rect 248607 11147 248641 11175
rect 248669 11147 248703 11175
rect 248731 11147 263877 11175
rect 263905 11147 263939 11175
rect 263967 11147 264001 11175
rect 264029 11147 264063 11175
rect 264091 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298990 11175
rect -958 11113 298990 11147
rect -958 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 171717 11113
rect 171745 11085 171779 11113
rect 171807 11085 171841 11113
rect 171869 11085 171903 11113
rect 171931 11085 187077 11113
rect 187105 11085 187139 11113
rect 187167 11085 187201 11113
rect 187229 11085 187263 11113
rect 187291 11085 202437 11113
rect 202465 11085 202499 11113
rect 202527 11085 202561 11113
rect 202589 11085 202623 11113
rect 202651 11085 217797 11113
rect 217825 11085 217859 11113
rect 217887 11085 217921 11113
rect 217949 11085 217983 11113
rect 218011 11085 233157 11113
rect 233185 11085 233219 11113
rect 233247 11085 233281 11113
rect 233309 11085 233343 11113
rect 233371 11085 248517 11113
rect 248545 11085 248579 11113
rect 248607 11085 248641 11113
rect 248669 11085 248703 11113
rect 248731 11085 263877 11113
rect 263905 11085 263939 11113
rect 263967 11085 264001 11113
rect 264029 11085 264063 11113
rect 264091 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298990 11113
rect -958 11051 298990 11085
rect -958 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 171717 11051
rect 171745 11023 171779 11051
rect 171807 11023 171841 11051
rect 171869 11023 171903 11051
rect 171931 11023 187077 11051
rect 187105 11023 187139 11051
rect 187167 11023 187201 11051
rect 187229 11023 187263 11051
rect 187291 11023 202437 11051
rect 202465 11023 202499 11051
rect 202527 11023 202561 11051
rect 202589 11023 202623 11051
rect 202651 11023 217797 11051
rect 217825 11023 217859 11051
rect 217887 11023 217921 11051
rect 217949 11023 217983 11051
rect 218011 11023 233157 11051
rect 233185 11023 233219 11051
rect 233247 11023 233281 11051
rect 233309 11023 233343 11051
rect 233371 11023 248517 11051
rect 248545 11023 248579 11051
rect 248607 11023 248641 11051
rect 248669 11023 248703 11051
rect 248731 11023 263877 11051
rect 263905 11023 263939 11051
rect 263967 11023 264001 11051
rect 264029 11023 264063 11051
rect 264091 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298990 11051
rect -958 10989 298990 11023
rect -958 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 171717 10989
rect 171745 10961 171779 10989
rect 171807 10961 171841 10989
rect 171869 10961 171903 10989
rect 171931 10961 187077 10989
rect 187105 10961 187139 10989
rect 187167 10961 187201 10989
rect 187229 10961 187263 10989
rect 187291 10961 202437 10989
rect 202465 10961 202499 10989
rect 202527 10961 202561 10989
rect 202589 10961 202623 10989
rect 202651 10961 217797 10989
rect 217825 10961 217859 10989
rect 217887 10961 217921 10989
rect 217949 10961 217983 10989
rect 218011 10961 233157 10989
rect 233185 10961 233219 10989
rect 233247 10961 233281 10989
rect 233309 10961 233343 10989
rect 233371 10961 248517 10989
rect 248545 10961 248579 10989
rect 248607 10961 248641 10989
rect 248669 10961 248703 10989
rect 248731 10961 263877 10989
rect 263905 10961 263939 10989
rect 263967 10961 264001 10989
rect 264029 10961 264063 10989
rect 264091 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298990 10989
rect -958 10913 298990 10961
rect -958 5175 298990 5223
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect -958 5113 298990 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect -958 5051 298990 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect -958 4989 298990 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect -958 4913 298990 4961
rect -958 2175 298990 2223
rect -958 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298990 2175
rect -958 2113 298990 2147
rect -958 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298990 2113
rect -958 2051 298990 2085
rect -958 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298990 2051
rect -958 1989 298990 2023
rect -958 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298990 1989
rect -958 1913 298990 1961
rect -478 -80 298510 -32
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect -478 -142 298510 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect -478 -204 298510 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect -478 -266 298510 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect -478 -342 298510 -294
rect -958 -560 298990 -512
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect -958 -622 298990 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect -958 -684 298990 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect -958 -746 298990 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect -958 -822 298990 -774
use user_proj_example  mprj
timestamp 0
transform 1 0 100000 0 1 100000
box 0 0 180000 178463
<< labels >>
flabel metal3 s 297780 3556 298500 3668 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 297780 201796 298500 201908 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 297780 221620 298500 221732 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 297780 241444 298500 241556 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 297780 261268 298500 261380 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 297780 281092 298500 281204 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 292348 297780 292460 298500 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 259252 297780 259364 298500 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 226156 297780 226268 298500 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 193060 297780 193172 298500 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 159964 297780 160076 298500 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 297780 23380 298500 23492 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 126868 297780 126980 298500 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 93772 297780 93884 298500 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 60676 297780 60788 298500 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 27580 297780 27692 298500 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -480 293580 240 293692 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -480 272412 240 272524 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -480 251244 240 251356 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -480 230076 240 230188 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -480 208908 240 209020 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -480 187740 240 187852 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 297780 43204 298500 43316 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -480 166572 240 166684 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -480 145404 240 145516 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -480 124236 240 124348 0 FreeSans 448 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -480 103068 240 103180 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -480 81900 240 82012 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -480 60732 240 60844 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -480 39564 240 39676 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -480 18396 240 18508 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 297780 63028 298500 63140 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 297780 82852 298500 82964 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 297780 102676 298500 102788 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 297780 122500 298500 122612 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 297780 142324 298500 142436 0 FreeSans 448 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 297780 162148 298500 162260 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 297780 181972 298500 182084 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 297780 16772 298500 16884 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 297780 215012 298500 215124 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 297780 234836 298500 234948 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 297780 254660 298500 254772 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 297780 274484 298500 274596 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 297780 294308 298500 294420 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 270284 297780 270396 298500 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 237188 297780 237300 298500 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 204092 297780 204204 298500 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 170996 297780 171108 298500 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 137900 297780 138012 298500 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 297780 36596 298500 36708 0 FreeSans 448 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 104804 297780 104916 298500 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 71708 297780 71820 298500 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 38612 297780 38724 298500 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 5516 297780 5628 298500 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -480 279468 240 279580 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -480 258300 240 258412 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -480 237132 240 237244 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -480 215964 240 216076 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -480 194796 240 194908 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -480 173628 240 173740 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 297780 56420 298500 56532 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -480 152460 240 152572 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -480 131292 240 131404 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -480 110124 240 110236 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -480 88956 240 89068 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -480 67788 240 67900 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -480 46620 240 46732 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -480 25452 240 25564 0 FreeSans 448 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -480 4284 240 4396 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 297780 76244 298500 76356 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 297780 96068 298500 96180 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 297780 115892 298500 116004 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 297780 135716 298500 135828 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 297780 155540 298500 155652 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 297780 175364 298500 175476 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 297780 195188 298500 195300 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 297780 10164 298500 10276 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 297780 208404 298500 208516 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 297780 228228 298500 228340 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 297780 248052 298500 248164 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 297780 267876 298500 267988 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 297780 287700 298500 287812 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 281316 297780 281428 298500 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 248220 297780 248332 298500 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 215124 297780 215236 298500 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 182028 297780 182140 298500 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 148932 297780 149044 298500 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 297780 29988 298500 30100 0 FreeSans 448 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 115836 297780 115948 298500 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 82740 297780 82852 298500 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 49644 297780 49756 298500 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 16548 297780 16660 298500 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -480 286524 240 286636 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -480 265356 240 265468 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -480 244188 240 244300 0 FreeSans 448 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -480 223020 240 223132 0 FreeSans 448 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -480 201852 240 201964 0 FreeSans 448 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -480 180684 240 180796 0 FreeSans 448 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 297780 49812 298500 49924 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -480 159516 240 159628 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -480 138348 240 138460 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -480 117180 240 117292 0 FreeSans 448 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -480 96012 240 96124 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -480 74844 240 74956 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -480 53676 240 53788 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -480 32508 240 32620 0 FreeSans 448 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -480 11340 240 11452 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 297780 69636 298500 69748 0 FreeSans 448 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 297780 89460 298500 89572 0 FreeSans 448 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 297780 109284 298500 109396 0 FreeSans 448 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 297780 129108 298500 129220 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 297780 148932 298500 149044 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 297780 168756 298500 168868 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 297780 188580 298500 188692 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 106596 -480 106708 240 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 135156 -480 135268 240 0 FreeSans 448 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 138012 -480 138124 240 0 FreeSans 448 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 140868 -480 140980 240 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 143724 -480 143836 240 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 146580 -480 146692 240 0 FreeSans 448 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 149436 -480 149548 240 0 FreeSans 448 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 152292 -480 152404 240 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 155148 -480 155260 240 0 FreeSans 448 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 158004 -480 158116 240 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 160860 -480 160972 240 0 FreeSans 448 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 109452 -480 109564 240 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 163716 -480 163828 240 0 FreeSans 448 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 166572 -480 166684 240 0 FreeSans 448 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 169428 -480 169540 240 0 FreeSans 448 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 172284 -480 172396 240 0 FreeSans 448 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 175140 -480 175252 240 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 177996 -480 178108 240 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 180852 -480 180964 240 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 183708 -480 183820 240 0 FreeSans 448 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 186564 -480 186676 240 0 FreeSans 448 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 189420 -480 189532 240 0 FreeSans 448 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 112308 -480 112420 240 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 192276 -480 192388 240 0 FreeSans 448 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 195132 -480 195244 240 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 197988 -480 198100 240 0 FreeSans 448 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 200844 -480 200956 240 0 FreeSans 448 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 203700 -480 203812 240 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 206556 -480 206668 240 0 FreeSans 448 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 209412 -480 209524 240 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 212268 -480 212380 240 0 FreeSans 448 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 215124 -480 215236 240 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 217980 -480 218092 240 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 115164 -480 115276 240 0 FreeSans 448 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 220836 -480 220948 240 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 223692 -480 223804 240 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 226548 -480 226660 240 0 FreeSans 448 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 229404 -480 229516 240 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 232260 -480 232372 240 0 FreeSans 448 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 235116 -480 235228 240 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 237972 -480 238084 240 0 FreeSans 448 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 240828 -480 240940 240 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 243684 -480 243796 240 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 246540 -480 246652 240 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 118020 -480 118132 240 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 249396 -480 249508 240 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 252252 -480 252364 240 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 255108 -480 255220 240 0 FreeSans 448 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 257964 -480 258076 240 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 260820 -480 260932 240 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 263676 -480 263788 240 0 FreeSans 448 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 266532 -480 266644 240 0 FreeSans 448 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 269388 -480 269500 240 0 FreeSans 448 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 272244 -480 272356 240 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 275100 -480 275212 240 0 FreeSans 448 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 120876 -480 120988 240 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 277956 -480 278068 240 0 FreeSans 448 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 280812 -480 280924 240 0 FreeSans 448 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 283668 -480 283780 240 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 286524 -480 286636 240 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 123732 -480 123844 240 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 126588 -480 126700 240 0 FreeSans 448 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 129444 -480 129556 240 0 FreeSans 448 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 132300 -480 132412 240 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 107548 -480 107660 240 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 136108 -480 136220 240 0 FreeSans 448 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 138964 -480 139076 240 0 FreeSans 448 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 141820 -480 141932 240 0 FreeSans 448 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 144676 -480 144788 240 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 147532 -480 147644 240 0 FreeSans 448 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 150388 -480 150500 240 0 FreeSans 448 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 153244 -480 153356 240 0 FreeSans 448 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 156100 -480 156212 240 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 158956 -480 159068 240 0 FreeSans 448 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 161812 -480 161924 240 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 110404 -480 110516 240 0 FreeSans 448 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 164668 -480 164780 240 0 FreeSans 448 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 167524 -480 167636 240 0 FreeSans 448 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 170380 -480 170492 240 0 FreeSans 448 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 173236 -480 173348 240 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 176092 -480 176204 240 0 FreeSans 448 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 178948 -480 179060 240 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 181804 -480 181916 240 0 FreeSans 448 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 184660 -480 184772 240 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 187516 -480 187628 240 0 FreeSans 448 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 190372 -480 190484 240 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 113260 -480 113372 240 0 FreeSans 448 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 193228 -480 193340 240 0 FreeSans 448 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 196084 -480 196196 240 0 FreeSans 448 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 198940 -480 199052 240 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 201796 -480 201908 240 0 FreeSans 448 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 204652 -480 204764 240 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 207508 -480 207620 240 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 210364 -480 210476 240 0 FreeSans 448 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 213220 -480 213332 240 0 FreeSans 448 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 216076 -480 216188 240 0 FreeSans 448 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 218932 -480 219044 240 0 FreeSans 448 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 116116 -480 116228 240 0 FreeSans 448 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 221788 -480 221900 240 0 FreeSans 448 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 224644 -480 224756 240 0 FreeSans 448 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 227500 -480 227612 240 0 FreeSans 448 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 230356 -480 230468 240 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 233212 -480 233324 240 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 236068 -480 236180 240 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 238924 -480 239036 240 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 241780 -480 241892 240 0 FreeSans 448 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 244636 -480 244748 240 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 247492 -480 247604 240 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 118972 -480 119084 240 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 250348 -480 250460 240 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 253204 -480 253316 240 0 FreeSans 448 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 256060 -480 256172 240 0 FreeSans 448 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 258916 -480 259028 240 0 FreeSans 448 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 261772 -480 261884 240 0 FreeSans 448 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 264628 -480 264740 240 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 267484 -480 267596 240 0 FreeSans 448 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 270340 -480 270452 240 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 273196 -480 273308 240 0 FreeSans 448 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 276052 -480 276164 240 0 FreeSans 448 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 121828 -480 121940 240 0 FreeSans 448 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 278908 -480 279020 240 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 281764 -480 281876 240 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 284620 -480 284732 240 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 287476 -480 287588 240 0 FreeSans 448 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 124684 -480 124796 240 0 FreeSans 448 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 127540 -480 127652 240 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 130396 -480 130508 240 0 FreeSans 448 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 133252 -480 133364 240 0 FreeSans 448 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 108500 -480 108612 240 0 FreeSans 448 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 137060 -480 137172 240 0 FreeSans 448 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 139916 -480 140028 240 0 FreeSans 448 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 142772 -480 142884 240 0 FreeSans 448 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 145628 -480 145740 240 0 FreeSans 448 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 148484 -480 148596 240 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 151340 -480 151452 240 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 154196 -480 154308 240 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 157052 -480 157164 240 0 FreeSans 448 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 159908 -480 160020 240 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 162764 -480 162876 240 0 FreeSans 448 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 111356 -480 111468 240 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 165620 -480 165732 240 0 FreeSans 448 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 168476 -480 168588 240 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 171332 -480 171444 240 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 174188 -480 174300 240 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 177044 -480 177156 240 0 FreeSans 448 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 179900 -480 180012 240 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 182756 -480 182868 240 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 185612 -480 185724 240 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 188468 -480 188580 240 0 FreeSans 448 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 191324 -480 191436 240 0 FreeSans 448 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 114212 -480 114324 240 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 194180 -480 194292 240 0 FreeSans 448 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 197036 -480 197148 240 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 199892 -480 200004 240 0 FreeSans 448 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 202748 -480 202860 240 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 205604 -480 205716 240 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 208460 -480 208572 240 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 211316 -480 211428 240 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 214172 -480 214284 240 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 217028 -480 217140 240 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 219884 -480 219996 240 0 FreeSans 448 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 117068 -480 117180 240 0 FreeSans 448 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 222740 -480 222852 240 0 FreeSans 448 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 225596 -480 225708 240 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 228452 -480 228564 240 0 FreeSans 448 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 231308 -480 231420 240 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 234164 -480 234276 240 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 237020 -480 237132 240 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 239876 -480 239988 240 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 242732 -480 242844 240 0 FreeSans 448 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 245588 -480 245700 240 0 FreeSans 448 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 248444 -480 248556 240 0 FreeSans 448 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 119924 -480 120036 240 0 FreeSans 448 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 251300 -480 251412 240 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 254156 -480 254268 240 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 257012 -480 257124 240 0 FreeSans 448 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 259868 -480 259980 240 0 FreeSans 448 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 262724 -480 262836 240 0 FreeSans 448 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 265580 -480 265692 240 0 FreeSans 448 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 268436 -480 268548 240 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 271292 -480 271404 240 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 274148 -480 274260 240 0 FreeSans 448 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 277004 -480 277116 240 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 122780 -480 122892 240 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 279860 -480 279972 240 0 FreeSans 448 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 282716 -480 282828 240 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 285572 -480 285684 240 0 FreeSans 448 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 288428 -480 288540 240 0 FreeSans 448 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 125636 -480 125748 240 0 FreeSans 448 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 128492 -480 128604 240 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 131348 -480 131460 240 0 FreeSans 448 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 134204 -480 134316 240 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 289380 -480 289492 240 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 290332 -480 290444 240 0 FreeSans 448 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 291284 -480 291396 240 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 292236 -480 292348 240 0 FreeSans 448 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -478 -342 -168 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 -342 298510 -32 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 298344 298510 298654 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 298200 -342 298510 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 2709 -822 3019 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 18069 -822 18379 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 33429 -822 33739 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 48789 -822 49099 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64149 -822 64459 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 79509 -822 79819 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 94869 -822 95179 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110229 -822 110539 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110229 276831 110539 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 125589 -822 125899 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 125589 276831 125899 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 140949 -822 141259 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 140949 276831 141259 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 156309 -822 156619 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 156309 276831 156619 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 171669 -822 171979 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 171669 276831 171979 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 -822 187339 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 276831 187339 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 202389 -822 202699 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 202389 276831 202699 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217749 -822 218059 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217749 276831 218059 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 233109 -822 233419 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 233109 276831 233419 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 -822 248779 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 276831 248779 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263829 -822 264139 100689 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263829 276831 264139 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 279189 -822 279499 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 294549 -822 294859 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 1913 298990 2223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 10913 298990 11223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 19913 298990 20223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 28913 298990 29223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 37913 298990 38223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 46913 298990 47223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 55913 298990 56223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 64913 298990 65223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 73913 298990 74223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 82913 298990 83223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 91913 298990 92223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 100913 298990 101223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 109913 298990 110223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 118913 298990 119223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 127913 298990 128223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 136913 298990 137223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 145913 298990 146223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 154913 298990 155223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 163913 298990 164223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 172913 298990 173223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 181913 298990 182223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 190913 298990 191223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 199913 298990 200223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 208913 298990 209223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 217913 298990 218223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 226913 298990 227223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 235913 298990 236223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 244913 298990 245223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 253913 298990 254223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 262913 298990 263223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 271913 298990 272223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 280913 298990 281223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 289913 298990 290223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -958 -822 -648 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 -822 298990 -512 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 298824 298990 299134 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 298680 -822 298990 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 4569 -822 4879 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 19929 -822 20239 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 35289 -822 35599 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50649 -822 50959 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66009 -822 66319 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 81369 -822 81679 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96729 -822 97039 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 -822 112399 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 276831 112399 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 127449 -822 127759 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 127449 276831 127759 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 142809 -822 143119 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 142809 276831 143119 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 158169 -822 158479 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 158169 276831 158479 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 -822 173839 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 276831 173839 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 -822 189199 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 276831 189199 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204249 -822 204559 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204249 276831 204559 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219609 -822 219919 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219609 276831 219919 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 234969 -822 235279 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 234969 276831 235279 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 -822 250639 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 276831 250639 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265689 -822 265999 100689 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265689 276831 265999 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 281049 -822 281359 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 296409 -822 296719 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 4913 298990 5223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 13913 298990 14223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 22913 298990 23223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 31913 298990 32223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 40913 298990 41223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 49913 298990 50223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 58913 298990 59223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 67913 298990 68223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 76913 298990 77223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 85913 298990 86223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 94913 298990 95223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 103913 298990 104223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 112913 298990 113223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 121913 298990 122223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 130913 298990 131223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 139913 298990 140223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 148913 298990 149223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 157913 298990 158223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 166913 298990 167223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 175913 298990 176223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 184913 298990 185223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 193913 298990 194223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 202913 298990 203223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 211913 298990 212223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 220913 298990 221223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 229913 298990 230223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 238913 298990 239223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 247913 298990 248223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 256913 298990 257223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 265913 298990 266223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 274913 298990 275223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 283913 298990 284223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 292913 298990 293223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 5684 -480 5796 240 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6636 -480 6748 240 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 7588 -480 7700 240 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 11396 -480 11508 240 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 43764 -480 43876 240 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 46620 -480 46732 240 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 49476 -480 49588 240 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 52332 -480 52444 240 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 55188 -480 55300 240 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 58044 -480 58156 240 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 60900 -480 61012 240 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 63756 -480 63868 240 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 66612 -480 66724 240 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 69468 -480 69580 240 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 15204 -480 15316 240 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 72324 -480 72436 240 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 75180 -480 75292 240 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 78036 -480 78148 240 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 80892 -480 81004 240 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 83748 -480 83860 240 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 86604 -480 86716 240 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 89460 -480 89572 240 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 92316 -480 92428 240 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 95172 -480 95284 240 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 98028 -480 98140 240 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 19012 -480 19124 240 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 100884 -480 100996 240 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 103740 -480 103852 240 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 22820 -480 22932 240 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 26628 -480 26740 240 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 29484 -480 29596 240 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 32340 -480 32452 240 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 35196 -480 35308 240 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 38052 -480 38164 240 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 40908 -480 41020 240 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 8540 -480 8652 240 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 12348 -480 12460 240 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 44716 -480 44828 240 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 47572 -480 47684 240 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 50428 -480 50540 240 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 53284 -480 53396 240 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 56140 -480 56252 240 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 58996 -480 59108 240 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 61852 -480 61964 240 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 64708 -480 64820 240 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 67564 -480 67676 240 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 70420 -480 70532 240 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 16156 -480 16268 240 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 73276 -480 73388 240 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 76132 -480 76244 240 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 78988 -480 79100 240 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 81844 -480 81956 240 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 84700 -480 84812 240 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 87556 -480 87668 240 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 90412 -480 90524 240 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 93268 -480 93380 240 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 96124 -480 96236 240 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 98980 -480 99092 240 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 19964 -480 20076 240 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 101836 -480 101948 240 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 104692 -480 104804 240 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 23772 -480 23884 240 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 27580 -480 27692 240 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 30436 -480 30548 240 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 33292 -480 33404 240 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 36148 -480 36260 240 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 39004 -480 39116 240 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 41860 -480 41972 240 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 13300 -480 13412 240 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 45668 -480 45780 240 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 48524 -480 48636 240 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 51380 -480 51492 240 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 54236 -480 54348 240 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 57092 -480 57204 240 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 59948 -480 60060 240 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 62804 -480 62916 240 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 65660 -480 65772 240 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 68516 -480 68628 240 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 71372 -480 71484 240 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 17108 -480 17220 240 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 74228 -480 74340 240 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 77084 -480 77196 240 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 79940 -480 80052 240 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 82796 -480 82908 240 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 85652 -480 85764 240 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 88508 -480 88620 240 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 91364 -480 91476 240 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 94220 -480 94332 240 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 97076 -480 97188 240 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 99932 -480 100044 240 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 20916 -480 21028 240 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 102788 -480 102900 240 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 105644 -480 105756 240 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 24724 -480 24836 240 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 28532 -480 28644 240 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 31388 -480 31500 240 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 34244 -480 34356 240 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 37100 -480 37212 240 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 39956 -480 40068 240 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 42812 -480 42924 240 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 14252 -480 14364 240 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 18060 -480 18172 240 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 21868 -480 21980 240 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 25676 -480 25788 240 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 9492 -480 9604 240 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 10444 -480 10556 240 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 279437 272161 279437 272161 0 vdd
rlabel via4 278975 275161 278975 275161 0 vss
rlabel metal4 281764 54264 281764 54264 0 io_in[0]
rlabel metal4 281876 75264 281876 75264 0 io_in[1]
rlabel metal4 282156 96264 282156 96264 0 io_in[2]
rlabel metal3 49455 166572 49455 166572 0 io_in[30]
rlabel metal3 49539 145404 49539 145404 0 io_in[31]
rlabel metal3 49511 124236 49511 124236 0 io_in[32]
rlabel metal3 49567 103068 49567 103068 0 io_in[33]
rlabel metal3 49427 81900 49427 81900 0 io_in[34]
rlabel metal3 49455 60732 49455 60732 0 io_in[35]
rlabel metal3 99449 141932 99449 141932 0 io_in[36]
rlabel metal3 99421 119756 99421 119756 0 io_in[37]
rlabel metal4 281988 117264 281988 117264 0 io_in[3]
rlabel metal3 281904 104916 281904 104916 0 io_in[4]
rlabel metal3 281848 119308 281848 119308 0 io_in[5]
rlabel metal2 281484 124684 281484 124684 0 io_in[6]
rlabel metal4 281876 201264 281876 201264 0 io_in[7]
rlabel metal4 282212 68292 282212 68292 0 io_oeb[0]
rlabel metal4 281820 89264 281820 89264 0 io_oeb[1]
rlabel metal4 282044 110264 282044 110264 0 io_oeb[2]
rlabel metal3 49483 152460 49483 152460 0 io_oeb[30]
rlabel metal3 49455 131292 49455 131292 0 io_oeb[31]
rlabel metal3 99505 215852 99505 215852 0 io_oeb[32]
rlabel metal3 49623 88956 49623 88956 0 io_oeb[33]
rlabel metal3 49651 67788 49651 67788 0 io_oeb[34]
rlabel metal3 49483 46620 49483 46620 0 io_oeb[35]
rlabel metal3 1267 25564 1267 25564 0 io_oeb[36]
rlabel metal3 1295 4396 1295 4396 0 io_oeb[37]
rlabel metal4 281932 131264 281932 131264 0 io_oeb[3]
rlabel metal4 282660 152264 282660 152264 0 io_oeb[4]
rlabel metal4 283500 173292 283500 173292 0 io_oeb[5]
rlabel metal4 284340 194264 284340 194264 0 io_oeb[6]
rlabel metal2 281428 155932 281428 155932 0 io_oeb[7]
rlabel metal4 285180 61264 285180 61264 0 io_out[0]
rlabel metal3 292761 29988 292761 29988 0 io_out[1]
rlabel metal4 282100 103264 282100 103264 0 io_out[2]
rlabel metal3 1155 159572 1155 159572 0 io_out[30]
rlabel metal3 1183 138460 1183 138460 0 io_out[31]
rlabel metal3 1211 117292 1211 117292 0 io_out[32]
rlabel metal3 1995 96124 1995 96124 0 io_out[33]
rlabel metal3 1239 74956 1239 74956 0 io_out[34]
rlabel metal3 1155 53732 1155 53732 0 io_out[35]
rlabel metal3 1183 32620 1183 32620 0 io_out[36]
rlabel metal3 1211 11452 1211 11452 0 io_out[37]
rlabel metal3 293601 69636 293601 69636 0 io_out[3]
rlabel metal3 295281 89572 295281 89572 0 io_out[4]
rlabel metal4 286020 166264 286020 166264 0 io_out[5]
rlabel metal3 292341 129108 292341 129108 0 io_out[6]
rlabel metal4 281820 208264 281820 208264 0 io_out[7]
rlabel metal3 106204 2548 106204 2548 0 la_data_in[0]
rlabel metal2 165956 51352 165956 51352 0 la_data_in[10]
rlabel metal2 138012 4095 138012 4095 0 la_data_in[11]
rlabel metal2 140980 1575 140980 1575 0 la_data_in[12]
rlabel metal2 143724 32235 143724 32235 0 la_data_in[13]
rlabel metal3 188300 98700 188300 98700 0 la_data_in[14]
rlabel metal2 190540 54873 190540 54873 0 la_data_in[15]
rlabel metal2 152292 3703 152292 3703 0 la_data_in[16]
rlabel metal2 155148 4515 155148 4515 0 la_data_in[17]
rlabel metal2 158116 1379 158116 1379 0 la_data_in[18]
rlabel metal3 179060 12180 179060 12180 0 la_data_in[19]
rlabel metal2 109452 6643 109452 6643 0 la_data_in[1]
rlabel metal2 163772 1631 163772 1631 0 la_data_in[20]
rlabel metal2 166572 6671 166572 6671 0 la_data_in[21]
rlabel metal2 202300 58205 202300 58205 0 la_data_in[22]
rlabel metal2 203980 57365 203980 57365 0 la_data_in[23]
rlabel metal2 175140 3255 175140 3255 0 la_data_in[24]
rlabel metal2 177996 38115 177996 38115 0 la_data_in[25]
rlabel metal3 194936 15596 194936 15596 0 la_data_in[26]
rlabel metal2 210700 54061 210700 54061 0 la_data_in[27]
rlabel metal2 186676 1379 186676 1379 0 la_data_in[28]
rlabel metal2 189532 1659 189532 1659 0 la_data_in[29]
rlabel metal2 168700 51905 168700 51905 0 la_data_in[2]
rlabel metal2 192332 1575 192332 1575 0 la_data_in[30]
rlabel metal3 212940 2940 212940 2940 0 la_data_in[31]
rlabel metal2 197988 3675 197988 3675 0 la_data_in[32]
rlabel metal2 200844 21315 200844 21315 0 la_data_in[33]
rlabel metal2 203700 4515 203700 4515 0 la_data_in[34]
rlabel metal2 224140 51541 224140 51541 0 la_data_in[35]
rlabel metal2 225820 51933 225820 51933 0 la_data_in[36]
rlabel metal2 212268 3255 212268 3255 0 la_data_in[37]
rlabel metal2 215236 1575 215236 1575 0 la_data_in[38]
rlabel metal2 218092 1575 218092 1575 0 la_data_in[39]
rlabel metal3 142772 14700 142772 14700 0 la_data_in[3]
rlabel metal2 220836 3675 220836 3675 0 la_data_in[40]
rlabel metal2 223804 1995 223804 1995 0 la_data_in[41]
rlabel metal2 226548 49035 226548 49035 0 la_data_in[42]
rlabel metal2 237580 51513 237580 51513 0 la_data_in[43]
rlabel metal2 239260 53165 239260 53165 0 la_data_in[44]
rlabel metal2 235172 1575 235172 1575 0 la_data_in[45]
rlabel metal2 238084 1295 238084 1295 0 la_data_in[46]
rlabel metal3 242564 99092 242564 99092 0 la_data_in[47]
rlabel metal2 245980 99197 245980 99197 0 la_data_in[48]
rlabel metal3 247128 99036 247128 99036 0 la_data_in[49]
rlabel metal2 118020 6223 118020 6223 0 la_data_in[4]
rlabel metal2 249368 10080 249368 10080 0 la_data_in[50]
rlabel metal2 251020 99197 251020 99197 0 la_data_in[51]
rlabel metal3 253904 2156 253904 2156 0 la_data_in[52]
rlabel metal2 257964 1351 257964 1351 0 la_data_in[53]
rlabel metal2 260820 1575 260820 1575 0 la_data_in[54]
rlabel metal3 258048 99092 258048 99092 0 la_data_in[55]
rlabel metal2 259420 53165 259420 53165 0 la_data_in[56]
rlabel metal2 269388 1603 269388 1603 0 la_data_in[57]
rlabel metal3 271180 2548 271180 2548 0 la_data_in[58]
rlabel metal3 270256 97916 270256 97916 0 la_data_in[59]
rlabel metal2 120876 7903 120876 7903 0 la_data_in[5]
rlabel metal2 266140 99365 266140 99365 0 la_data_in[60]
rlabel metal2 280812 1603 280812 1603 0 la_data_in[61]
rlabel metal2 269500 98525 269500 98525 0 la_data_in[62]
rlabel metal2 271180 98945 271180 98945 0 la_data_in[63]
rlabel metal2 175420 58625 175420 58625 0 la_data_in[6]
rlabel metal2 177100 59073 177100 59073 0 la_data_in[7]
rlabel metal2 129444 9583 129444 9583 0 la_data_in[8]
rlabel metal2 132356 10843 132356 10843 0 la_data_in[9]
rlabel metal2 107548 4935 107548 4935 0 la_data_out[0]
rlabel metal2 136108 3675 136108 3675 0 la_data_out[10]
rlabel metal3 161672 22316 161672 22316 0 la_data_out[11]
rlabel metal2 141932 1631 141932 1631 0 la_data_out[12]
rlabel metal2 144676 4599 144676 4599 0 la_data_out[13]
rlabel metal2 189420 98945 189420 98945 0 la_data_out[14]
rlabel metal2 191100 62013 191100 62013 0 la_data_out[15]
rlabel metal2 153244 4123 153244 4123 0 la_data_out[16]
rlabel metal2 156100 12523 156100 12523 0 la_data_out[17]
rlabel metal2 158956 3311 158956 3311 0 la_data_out[18]
rlabel metal2 161812 4991 161812 4991 0 la_data_out[19]
rlabel metal2 167580 52381 167580 52381 0 la_data_out[1]
rlabel metal2 164780 2443 164780 2443 0 la_data_out[20]
rlabel metal2 167636 2051 167636 2051 0 la_data_out[21]
rlabel metal3 200760 99092 200760 99092 0 la_data_out[22]
rlabel metal2 173348 1995 173348 1995 0 la_data_out[23]
rlabel metal2 176204 2023 176204 2023 0 la_data_out[24]
rlabel metal2 178948 9135 178948 9135 0 la_data_out[25]
rlabel metal2 181804 3731 181804 3731 0 la_data_out[26]
rlabel metal2 211260 54453 211260 54453 0 la_data_out[27]
rlabel metal2 187516 4935 187516 4935 0 la_data_out[28]
rlabel metal2 190372 3283 190372 3283 0 la_data_out[29]
rlabel metal2 113316 8295 113316 8295 0 la_data_out[2]
rlabel metal2 193228 4123 193228 4123 0 la_data_out[30]
rlabel metal2 196084 9555 196084 9555 0 la_data_out[31]
rlabel metal2 198940 6195 198940 6195 0 la_data_out[32]
rlabel metal2 201796 6615 201796 6615 0 la_data_out[33]
rlabel metal2 223020 99169 223020 99169 0 la_data_out[34]
rlabel metal2 224700 54005 224700 54005 0 la_data_out[35]
rlabel metal2 210364 4963 210364 4963 0 la_data_out[36]
rlabel metal2 213220 6223 213220 6223 0 la_data_out[37]
rlabel metal2 216188 2415 216188 2415 0 la_data_out[38]
rlabel metal2 218932 3283 218932 3283 0 la_data_out[39]
rlabel metal2 116116 12915 116116 12915 0 la_data_out[3]
rlabel metal2 221900 1603 221900 1603 0 la_data_out[40]
rlabel metal2 224644 48615 224644 48615 0 la_data_out[41]
rlabel metal2 227612 1183 227612 1183 0 la_data_out[42]
rlabel metal2 238140 51121 238140 51121 0 la_data_out[43]
rlabel metal2 233324 1267 233324 1267 0 la_data_out[44]
rlabel metal2 236180 1155 236180 1155 0 la_data_out[45]
rlabel metal2 239036 1211 239036 1211 0 la_data_out[46]
rlabel metal2 241892 1155 241892 1155 0 la_data_out[47]
rlabel metal2 246540 99169 246540 99169 0 la_data_out[48]
rlabel metal3 247856 99092 247856 99092 0 la_data_out[49]
rlabel metal2 118972 13335 118972 13335 0 la_data_out[4]
rlabel metal3 250124 2100 250124 2100 0 la_data_out[50]
rlabel metal3 252392 99092 252392 99092 0 la_data_out[51]
rlabel metal2 256032 92400 256032 92400 0 la_data_out[52]
rlabel metal2 258916 1155 258916 1155 0 la_data_out[53]
rlabel metal2 261772 49455 261772 49455 0 la_data_out[54]
rlabel metal2 258300 75845 258300 75845 0 la_data_out[55]
rlabel metal2 259980 53585 259980 53585 0 la_data_out[56]
rlabel metal2 270340 2023 270340 2023 0 la_data_out[57]
rlabel metal2 273196 1995 273196 1995 0 la_data_out[58]
rlabel metal2 265020 54005 265020 54005 0 la_data_out[59]
rlabel metal3 148064 27300 148064 27300 0 la_data_out[5]
rlabel metal2 278908 1575 278908 1575 0 la_data_out[60]
rlabel metal2 281764 3255 281764 3255 0 la_data_out[61]
rlabel metal2 270060 98105 270060 98105 0 la_data_out[62]
rlabel metal2 271740 53585 271740 53585 0 la_data_out[63]
rlabel metal2 175980 55265 175980 55265 0 la_data_out[6]
rlabel metal2 177660 99505 177660 99505 0 la_data_out[7]
rlabel metal2 130396 14175 130396 14175 0 la_data_out[8]
rlabel metal2 133252 7875 133252 7875 0 la_data_out[9]
rlabel metal2 108500 15015 108500 15015 0 la_oenb[0]
rlabel metal2 177660 64792 177660 64792 0 la_oenb[10]
rlabel metal2 140028 2835 140028 2835 0 la_oenb[11]
rlabel metal2 142884 1603 142884 1603 0 la_oenb[12]
rlabel metal2 188300 56525 188300 56525 0 la_oenb[13]
rlabel metal2 189980 57393 189980 57393 0 la_oenb[14]
rlabel metal2 151340 9555 151340 9555 0 la_oenb[15]
rlabel metal2 154196 33103 154196 33103 0 la_oenb[16]
rlabel metal3 176064 25676 176064 25676 0 la_oenb[17]
rlabel metal3 177604 10556 177604 10556 0 la_oenb[18]
rlabel metal2 198380 84665 198380 84665 0 la_oenb[19]
rlabel metal2 168140 62405 168140 62405 0 la_oenb[1]
rlabel metal2 165620 6251 165620 6251 0 la_oenb[20]
rlabel metal2 168476 13363 168476 13363 0 la_oenb[21]
rlabel metal2 203420 63693 203420 63693 0 la_oenb[22]
rlabel metal2 174188 10815 174188 10815 0 la_oenb[23]
rlabel metal2 177044 8715 177044 8715 0 la_oenb[24]
rlabel metal2 180012 1155 180012 1155 0 la_oenb[25]
rlabel metal2 210140 64925 210140 64925 0 la_oenb[26]
rlabel metal2 211820 61145 211820 61145 0 la_oenb[27]
rlabel metal2 188580 1155 188580 1155 0 la_oenb[28]
rlabel metal2 191436 1351 191436 1351 0 la_oenb[29]
rlabel metal3 142044 23940 142044 23940 0 la_oenb[2]
rlabel metal2 194292 1155 194292 1155 0 la_oenb[30]
rlabel metal3 207788 25620 207788 25620 0 la_oenb[31]
rlabel metal2 199948 5355 199948 5355 0 la_oenb[32]
rlabel metal2 202860 1155 202860 1155 0 la_oenb[33]
rlabel metal2 223580 60725 223580 60725 0 la_oenb[34]
rlabel metal2 225260 51065 225260 51065 0 la_oenb[35]
rlabel metal2 211428 1183 211428 1183 0 la_oenb[36]
rlabel metal2 214284 1211 214284 1211 0 la_oenb[37]
rlabel metal2 217140 1239 217140 1239 0 la_oenb[38]
rlabel metal2 219996 1267 219996 1267 0 la_oenb[39]
rlabel metal2 117068 48615 117068 48615 0 la_oenb[3]
rlabel metal2 222740 49483 222740 49483 0 la_oenb[40]
rlabel metal2 225708 1155 225708 1155 0 la_oenb[41]
rlabel metal2 237020 99421 237020 99421 0 la_oenb[42]
rlabel metal2 238700 51149 238700 51149 0 la_oenb[43]
rlabel metal2 234164 49455 234164 49455 0 la_oenb[44]
rlabel metal2 237132 1183 237132 1183 0 la_oenb[45]
rlabel metal3 241808 99036 241808 99036 0 la_oenb[46]
rlabel metal2 245420 51261 245420 51261 0 la_oenb[47]
rlabel metal3 246344 99092 246344 99092 0 la_oenb[48]
rlabel metal2 248444 49245 248444 49245 0 la_oenb[49]
rlabel metal2 119924 8743 119924 8743 0 la_oenb[4]
rlabel metal2 250460 99169 250460 99169 0 la_oenb[50]
rlabel metal3 253148 99036 253148 99036 0 la_oenb[51]
rlabel metal2 257068 49315 257068 49315 0 la_oenb[52]
rlabel metal2 259868 49483 259868 49483 0 la_oenb[53]
rlabel metal3 259952 2044 259952 2044 0 la_oenb[54]
rlabel metal2 258860 51093 258860 51093 0 la_oenb[55]
rlabel metal2 260540 51065 260540 51065 0 la_oenb[56]
rlabel metal2 262220 60725 262220 60725 0 la_oenb[57]
rlabel metal2 274148 25935 274148 25935 0 la_oenb[58]
rlabel metal3 271880 93660 271880 93660 0 la_oenb[59]
rlabel metal2 174860 51933 174860 51933 0 la_oenb[5]
rlabel metal3 273560 27300 273560 27300 0 la_oenb[60]
rlabel metal2 268940 72065 268940 72065 0 la_oenb[61]
rlabel metal2 285628 1267 285628 1267 0 la_oenb[62]
rlabel metal2 272300 51149 272300 51149 0 la_oenb[63]
rlabel metal3 176288 99092 176288 99092 0 la_oenb[6]
rlabel metal2 128548 17143 128548 17143 0 la_oenb[7]
rlabel metal2 131348 8323 131348 8323 0 la_oenb[8]
rlabel metal2 134204 16695 134204 16695 0 la_oenb[9]
rlabel metal2 272860 51121 272860 51121 0 user_irq[0]
rlabel metal2 273420 51093 273420 51093 0 user_irq[1]
rlabel metal2 273980 51065 273980 51065 0 user_irq[2]
rlabel metal2 105980 99365 105980 99365 0 wb_clk_i
rlabel metal2 106540 63665 106540 63665 0 wb_rst_i
rlabel metal2 107100 54845 107100 54845 0 wbs_ack_o
rlabel metal2 11396 49035 11396 49035 0 wbs_adr_i[0]
rlabel metal2 128380 99169 128380 99169 0 wbs_adr_i[10]
rlabel metal2 46620 46935 46620 46935 0 wbs_adr_i[11]
rlabel metal2 49532 1603 49532 1603 0 wbs_adr_i[12]
rlabel metal2 133420 96425 133420 96425 0 wbs_adr_i[13]
rlabel metal2 55188 45675 55188 45675 0 wbs_adr_i[14]
rlabel metal2 58156 1575 58156 1575 0 wbs_adr_i[15]
rlabel metal2 61012 1603 61012 1603 0 wbs_adr_i[16]
rlabel metal2 140140 51541 140140 51541 0 wbs_adr_i[17]
rlabel metal2 141820 99505 141820 99505 0 wbs_adr_i[18]
rlabel metal2 69468 44835 69468 44835 0 wbs_adr_i[19]
rlabel metal2 15204 48615 15204 48615 0 wbs_adr_i[1]
rlabel metal2 72324 43995 72324 43995 0 wbs_adr_i[20]
rlabel metal2 75180 43603 75180 43603 0 wbs_adr_i[21]
rlabel metal3 113288 85260 113288 85260 0 wbs_adr_i[22]
rlabel metal2 80892 6223 80892 6223 0 wbs_adr_i[23]
rlabel metal2 83748 42343 83748 42343 0 wbs_adr_i[24]
rlabel metal2 153580 98973 153580 98973 0 wbs_adr_i[25]
rlabel metal2 155260 94325 155260 94325 0 wbs_adr_i[26]
rlabel metal3 156408 99092 156408 99092 0 wbs_adr_i[27]
rlabel metal2 95284 1379 95284 1379 0 wbs_adr_i[28]
rlabel metal2 98028 48223 98028 48223 0 wbs_adr_i[29]
rlabel metal2 19012 27195 19012 27195 0 wbs_adr_i[2]
rlabel metal3 131432 81900 131432 81900 0 wbs_adr_i[30]
rlabel metal2 163660 96873 163660 96873 0 wbs_adr_i[31]
rlabel metal2 22820 40215 22820 40215 0 wbs_adr_i[3]
rlabel metal2 26628 39795 26628 39795 0 wbs_adr_i[4]
rlabel metal2 119980 89285 119980 89285 0 wbs_adr_i[5]
rlabel metal2 121660 88865 121660 88865 0 wbs_adr_i[6]
rlabel metal2 35196 38115 35196 38115 0 wbs_adr_i[7]
rlabel metal2 38052 37695 38052 37695 0 wbs_adr_i[8]
rlabel metal2 41020 2051 41020 2051 0 wbs_adr_i[9]
rlabel metal2 107660 51905 107660 51905 0 wbs_cyc_i
rlabel metal2 12460 2023 12460 2023 0 wbs_dat_i[0]
rlabel metal2 128940 67025 128940 67025 0 wbs_dat_i[10]
rlabel metal2 47572 27615 47572 27615 0 wbs_dat_i[11]
rlabel metal2 50428 6615 50428 6615 0 wbs_dat_i[12]
rlabel metal3 93632 34860 93632 34860 0 wbs_dat_i[13]
rlabel metal2 56140 28455 56140 28455 0 wbs_dat_i[14]
rlabel metal2 58996 15435 58996 15435 0 wbs_dat_i[15]
rlabel metal2 61852 22575 61852 22575 0 wbs_dat_i[16]
rlabel metal2 140700 99169 140700 99169 0 wbs_dat_i[17]
rlabel metal2 142380 78785 142380 78785 0 wbs_dat_i[18]
rlabel metal2 70420 3311 70420 3311 0 wbs_dat_i[19]
rlabel metal2 16268 2443 16268 2443 0 wbs_dat_i[1]
rlabel metal2 73276 36015 73276 36015 0 wbs_dat_i[20]
rlabel metal3 111776 70980 111776 70980 0 wbs_dat_i[21]
rlabel metal2 78988 4963 78988 4963 0 wbs_dat_i[22]
rlabel metal2 81844 9555 81844 9555 0 wbs_dat_i[23]
rlabel metal2 84700 3731 84700 3731 0 wbs_dat_i[24]
rlabel metal2 154140 82985 154140 82985 0 wbs_dat_i[25]
rlabel metal2 155820 68285 155820 68285 0 wbs_dat_i[26]
rlabel metal2 93268 25935 93268 25935 0 wbs_dat_i[27]
rlabel metal2 96124 11235 96124 11235 0 wbs_dat_i[28]
rlabel metal2 98980 9135 98980 9135 0 wbs_dat_i[29]
rlabel metal2 20076 1127 20076 1127 0 wbs_dat_i[2]
rlabel metal3 132188 69300 132188 69300 0 wbs_dat_i[30]
rlabel metal2 104692 17955 104692 17955 0 wbs_dat_i[31]
rlabel metal2 23772 26355 23772 26355 0 wbs_dat_i[3]
rlabel metal2 27580 13335 27580 13335 0 wbs_dat_i[4]
rlabel metal2 120540 66605 120540 66605 0 wbs_dat_i[5]
rlabel metal2 33404 2835 33404 2835 0 wbs_dat_i[6]
rlabel metal2 36148 3255 36148 3255 0 wbs_dat_i[7]
rlabel metal2 39004 3283 39004 3283 0 wbs_dat_i[8]
rlabel metal2 41860 3675 41860 3675 0 wbs_dat_i[9]
rlabel metal2 13412 2415 13412 2415 0 wbs_dat_o[0]
rlabel metal2 45668 3703 45668 3703 0 wbs_dat_o[10]
rlabel metal2 48524 21735 48524 21735 0 wbs_dat_o[11]
rlabel metal2 132860 79205 132860 79205 0 wbs_dat_o[12]
rlabel metal2 54236 4095 54236 4095 0 wbs_dat_o[13]
rlabel metal2 57148 4123 57148 4123 0 wbs_dat_o[14]
rlabel metal2 59948 4151 59948 4151 0 wbs_dat_o[15]
rlabel metal2 62804 35175 62804 35175 0 wbs_dat_o[16]
rlabel metal2 141260 99365 141260 99365 0 wbs_dat_o[17]
rlabel metal2 142772 97678 142772 97678 0 wbs_dat_o[18]
rlabel metal2 71428 4515 71428 4515 0 wbs_dat_o[19]
rlabel metal3 64904 84420 64904 84420 0 wbs_dat_o[1]
rlabel metal2 74228 4543 74228 4543 0 wbs_dat_o[20]
rlabel metal3 112532 37380 112532 37380 0 wbs_dat_o[21]
rlabel metal2 79940 4571 79940 4571 0 wbs_dat_o[22]
rlabel metal2 82796 26775 82796 26775 0 wbs_dat_o[23]
rlabel metal2 85708 22155 85708 22155 0 wbs_dat_o[24]
rlabel metal2 154700 80045 154700 80045 0 wbs_dat_o[25]
rlabel metal3 155288 99036 155288 99036 0 wbs_dat_o[26]
rlabel metal2 94220 45703 94220 45703 0 wbs_dat_o[27]
rlabel metal2 97188 735 97188 735 0 wbs_dat_o[28]
rlabel metal3 130704 39060 130704 39060 0 wbs_dat_o[29]
rlabel metal3 67928 14700 67928 14700 0 wbs_dat_o[2]
rlabel metal2 163100 69965 163100 69965 0 wbs_dat_o[30]
rlabel metal2 105644 10815 105644 10815 0 wbs_dat_o[31]
rlabel metal2 24724 43575 24724 43575 0 wbs_dat_o[3]
rlabel metal2 119420 64085 119420 64085 0 wbs_dat_o[4]
rlabel metal2 121100 71225 121100 71225 0 wbs_dat_o[5]
rlabel metal2 34244 7875 34244 7875 0 wbs_dat_o[6]
rlabel metal2 37100 24255 37100 24255 0 wbs_dat_o[7]
rlabel metal2 39956 33495 39956 33495 0 wbs_dat_o[8]
rlabel metal2 127820 82145 127820 82145 0 wbs_dat_o[9]
rlabel metal2 14308 30975 14308 30975 0 wbs_sel_i[0]
rlabel metal2 18172 1211 18172 1211 0 wbs_sel_i[1]
rlabel metal2 21980 1239 21980 1239 0 wbs_sel_i[2]
rlabel metal2 25788 1267 25788 1267 0 wbs_sel_i[3]
rlabel metal2 108220 51065 108220 51065 0 wbs_stb_i
rlabel metal2 10556 1183 10556 1183 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 298020 298020
<< end >>
