magic
tech gf180mcuD
magscale 1 5
timestamp 1701943170
<< obsm1 >>
rect 672 463 179312 178457
<< metal2 >>
rect 5936 0 5992 400
rect 6496 0 6552 400
rect 7056 0 7112 400
rect 7616 0 7672 400
rect 8176 0 8232 400
rect 8736 0 8792 400
rect 9296 0 9352 400
rect 9856 0 9912 400
rect 10416 0 10472 400
rect 10976 0 11032 400
rect 11536 0 11592 400
rect 12096 0 12152 400
rect 12656 0 12712 400
rect 13216 0 13272 400
rect 13776 0 13832 400
rect 14336 0 14392 400
rect 14896 0 14952 400
rect 15456 0 15512 400
rect 16016 0 16072 400
rect 16576 0 16632 400
rect 17136 0 17192 400
rect 17696 0 17752 400
rect 18256 0 18312 400
rect 18816 0 18872 400
rect 19376 0 19432 400
rect 19936 0 19992 400
rect 20496 0 20552 400
rect 21056 0 21112 400
rect 21616 0 21672 400
rect 22176 0 22232 400
rect 22736 0 22792 400
rect 23296 0 23352 400
rect 23856 0 23912 400
rect 24416 0 24472 400
rect 24976 0 25032 400
rect 25536 0 25592 400
rect 26096 0 26152 400
rect 26656 0 26712 400
rect 27216 0 27272 400
rect 27776 0 27832 400
rect 28336 0 28392 400
rect 28896 0 28952 400
rect 29456 0 29512 400
rect 30016 0 30072 400
rect 30576 0 30632 400
rect 31136 0 31192 400
rect 31696 0 31752 400
rect 32256 0 32312 400
rect 32816 0 32872 400
rect 33376 0 33432 400
rect 33936 0 33992 400
rect 34496 0 34552 400
rect 35056 0 35112 400
rect 35616 0 35672 400
rect 36176 0 36232 400
rect 36736 0 36792 400
rect 37296 0 37352 400
rect 37856 0 37912 400
rect 38416 0 38472 400
rect 38976 0 39032 400
rect 39536 0 39592 400
rect 40096 0 40152 400
rect 40656 0 40712 400
rect 41216 0 41272 400
rect 41776 0 41832 400
rect 42336 0 42392 400
rect 42896 0 42952 400
rect 43456 0 43512 400
rect 44016 0 44072 400
rect 44576 0 44632 400
rect 45136 0 45192 400
rect 45696 0 45752 400
rect 46256 0 46312 400
rect 46816 0 46872 400
rect 47376 0 47432 400
rect 47936 0 47992 400
rect 48496 0 48552 400
rect 49056 0 49112 400
rect 49616 0 49672 400
rect 50176 0 50232 400
rect 50736 0 50792 400
rect 51296 0 51352 400
rect 51856 0 51912 400
rect 52416 0 52472 400
rect 52976 0 53032 400
rect 53536 0 53592 400
rect 54096 0 54152 400
rect 54656 0 54712 400
rect 55216 0 55272 400
rect 55776 0 55832 400
rect 56336 0 56392 400
rect 56896 0 56952 400
rect 57456 0 57512 400
rect 58016 0 58072 400
rect 58576 0 58632 400
rect 59136 0 59192 400
rect 59696 0 59752 400
rect 60256 0 60312 400
rect 60816 0 60872 400
rect 61376 0 61432 400
rect 61936 0 61992 400
rect 62496 0 62552 400
rect 63056 0 63112 400
rect 63616 0 63672 400
rect 64176 0 64232 400
rect 64736 0 64792 400
rect 65296 0 65352 400
rect 65856 0 65912 400
rect 66416 0 66472 400
rect 66976 0 67032 400
rect 67536 0 67592 400
rect 68096 0 68152 400
rect 68656 0 68712 400
rect 69216 0 69272 400
rect 69776 0 69832 400
rect 70336 0 70392 400
rect 70896 0 70952 400
rect 71456 0 71512 400
rect 72016 0 72072 400
rect 72576 0 72632 400
rect 73136 0 73192 400
rect 73696 0 73752 400
rect 74256 0 74312 400
rect 74816 0 74872 400
rect 75376 0 75432 400
rect 75936 0 75992 400
rect 76496 0 76552 400
rect 77056 0 77112 400
rect 77616 0 77672 400
rect 78176 0 78232 400
rect 78736 0 78792 400
rect 79296 0 79352 400
rect 79856 0 79912 400
rect 80416 0 80472 400
rect 80976 0 81032 400
rect 81536 0 81592 400
rect 82096 0 82152 400
rect 82656 0 82712 400
rect 83216 0 83272 400
rect 83776 0 83832 400
rect 84336 0 84392 400
rect 84896 0 84952 400
rect 85456 0 85512 400
rect 86016 0 86072 400
rect 86576 0 86632 400
rect 87136 0 87192 400
rect 87696 0 87752 400
rect 88256 0 88312 400
rect 88816 0 88872 400
rect 89376 0 89432 400
rect 89936 0 89992 400
rect 90496 0 90552 400
rect 91056 0 91112 400
rect 91616 0 91672 400
rect 92176 0 92232 400
rect 92736 0 92792 400
rect 93296 0 93352 400
rect 93856 0 93912 400
rect 94416 0 94472 400
rect 94976 0 95032 400
rect 95536 0 95592 400
rect 96096 0 96152 400
rect 96656 0 96712 400
rect 97216 0 97272 400
rect 97776 0 97832 400
rect 98336 0 98392 400
rect 98896 0 98952 400
rect 99456 0 99512 400
rect 100016 0 100072 400
rect 100576 0 100632 400
rect 101136 0 101192 400
rect 101696 0 101752 400
rect 102256 0 102312 400
rect 102816 0 102872 400
rect 103376 0 103432 400
rect 103936 0 103992 400
rect 104496 0 104552 400
rect 105056 0 105112 400
rect 105616 0 105672 400
rect 106176 0 106232 400
rect 106736 0 106792 400
rect 107296 0 107352 400
rect 107856 0 107912 400
rect 108416 0 108472 400
rect 108976 0 109032 400
rect 109536 0 109592 400
rect 110096 0 110152 400
rect 110656 0 110712 400
rect 111216 0 111272 400
rect 111776 0 111832 400
rect 112336 0 112392 400
rect 112896 0 112952 400
rect 113456 0 113512 400
rect 114016 0 114072 400
rect 114576 0 114632 400
rect 115136 0 115192 400
rect 115696 0 115752 400
rect 116256 0 116312 400
rect 116816 0 116872 400
rect 117376 0 117432 400
rect 117936 0 117992 400
rect 118496 0 118552 400
rect 119056 0 119112 400
rect 119616 0 119672 400
rect 120176 0 120232 400
rect 120736 0 120792 400
rect 121296 0 121352 400
rect 121856 0 121912 400
rect 122416 0 122472 400
rect 122976 0 123032 400
rect 123536 0 123592 400
rect 124096 0 124152 400
rect 124656 0 124712 400
rect 125216 0 125272 400
rect 125776 0 125832 400
rect 126336 0 126392 400
rect 126896 0 126952 400
rect 127456 0 127512 400
rect 128016 0 128072 400
rect 128576 0 128632 400
rect 129136 0 129192 400
rect 129696 0 129752 400
rect 130256 0 130312 400
rect 130816 0 130872 400
rect 131376 0 131432 400
rect 131936 0 131992 400
rect 132496 0 132552 400
rect 133056 0 133112 400
rect 133616 0 133672 400
rect 134176 0 134232 400
rect 134736 0 134792 400
rect 135296 0 135352 400
rect 135856 0 135912 400
rect 136416 0 136472 400
rect 136976 0 137032 400
rect 137536 0 137592 400
rect 138096 0 138152 400
rect 138656 0 138712 400
rect 139216 0 139272 400
rect 139776 0 139832 400
rect 140336 0 140392 400
rect 140896 0 140952 400
rect 141456 0 141512 400
rect 142016 0 142072 400
rect 142576 0 142632 400
rect 143136 0 143192 400
rect 143696 0 143752 400
rect 144256 0 144312 400
rect 144816 0 144872 400
rect 145376 0 145432 400
rect 145936 0 145992 400
rect 146496 0 146552 400
rect 147056 0 147112 400
rect 147616 0 147672 400
rect 148176 0 148232 400
rect 148736 0 148792 400
rect 149296 0 149352 400
rect 149856 0 149912 400
rect 150416 0 150472 400
rect 150976 0 151032 400
rect 151536 0 151592 400
rect 152096 0 152152 400
rect 152656 0 152712 400
rect 153216 0 153272 400
rect 153776 0 153832 400
rect 154336 0 154392 400
rect 154896 0 154952 400
rect 155456 0 155512 400
rect 156016 0 156072 400
rect 156576 0 156632 400
rect 157136 0 157192 400
rect 157696 0 157752 400
rect 158256 0 158312 400
rect 158816 0 158872 400
rect 159376 0 159432 400
rect 159936 0 159992 400
rect 160496 0 160552 400
rect 161056 0 161112 400
rect 161616 0 161672 400
rect 162176 0 162232 400
rect 162736 0 162792 400
rect 163296 0 163352 400
rect 163856 0 163912 400
rect 164416 0 164472 400
rect 164976 0 165032 400
rect 165536 0 165592 400
rect 166096 0 166152 400
rect 166656 0 166712 400
rect 167216 0 167272 400
rect 167776 0 167832 400
rect 168336 0 168392 400
rect 168896 0 168952 400
rect 169456 0 169512 400
rect 170016 0 170072 400
rect 170576 0 170632 400
rect 171136 0 171192 400
rect 171696 0 171752 400
rect 172256 0 172312 400
rect 172816 0 172872 400
rect 173376 0 173432 400
rect 173936 0 173992 400
<< obsm2 >>
rect 630 430 179130 178463
rect 630 350 5906 430
rect 6022 350 6466 430
rect 6582 350 7026 430
rect 7142 350 7586 430
rect 7702 350 8146 430
rect 8262 350 8706 430
rect 8822 350 9266 430
rect 9382 350 9826 430
rect 9942 350 10386 430
rect 10502 350 10946 430
rect 11062 350 11506 430
rect 11622 350 12066 430
rect 12182 350 12626 430
rect 12742 350 13186 430
rect 13302 350 13746 430
rect 13862 350 14306 430
rect 14422 350 14866 430
rect 14982 350 15426 430
rect 15542 350 15986 430
rect 16102 350 16546 430
rect 16662 350 17106 430
rect 17222 350 17666 430
rect 17782 350 18226 430
rect 18342 350 18786 430
rect 18902 350 19346 430
rect 19462 350 19906 430
rect 20022 350 20466 430
rect 20582 350 21026 430
rect 21142 350 21586 430
rect 21702 350 22146 430
rect 22262 350 22706 430
rect 22822 350 23266 430
rect 23382 350 23826 430
rect 23942 350 24386 430
rect 24502 350 24946 430
rect 25062 350 25506 430
rect 25622 350 26066 430
rect 26182 350 26626 430
rect 26742 350 27186 430
rect 27302 350 27746 430
rect 27862 350 28306 430
rect 28422 350 28866 430
rect 28982 350 29426 430
rect 29542 350 29986 430
rect 30102 350 30546 430
rect 30662 350 31106 430
rect 31222 350 31666 430
rect 31782 350 32226 430
rect 32342 350 32786 430
rect 32902 350 33346 430
rect 33462 350 33906 430
rect 34022 350 34466 430
rect 34582 350 35026 430
rect 35142 350 35586 430
rect 35702 350 36146 430
rect 36262 350 36706 430
rect 36822 350 37266 430
rect 37382 350 37826 430
rect 37942 350 38386 430
rect 38502 350 38946 430
rect 39062 350 39506 430
rect 39622 350 40066 430
rect 40182 350 40626 430
rect 40742 350 41186 430
rect 41302 350 41746 430
rect 41862 350 42306 430
rect 42422 350 42866 430
rect 42982 350 43426 430
rect 43542 350 43986 430
rect 44102 350 44546 430
rect 44662 350 45106 430
rect 45222 350 45666 430
rect 45782 350 46226 430
rect 46342 350 46786 430
rect 46902 350 47346 430
rect 47462 350 47906 430
rect 48022 350 48466 430
rect 48582 350 49026 430
rect 49142 350 49586 430
rect 49702 350 50146 430
rect 50262 350 50706 430
rect 50822 350 51266 430
rect 51382 350 51826 430
rect 51942 350 52386 430
rect 52502 350 52946 430
rect 53062 350 53506 430
rect 53622 350 54066 430
rect 54182 350 54626 430
rect 54742 350 55186 430
rect 55302 350 55746 430
rect 55862 350 56306 430
rect 56422 350 56866 430
rect 56982 350 57426 430
rect 57542 350 57986 430
rect 58102 350 58546 430
rect 58662 350 59106 430
rect 59222 350 59666 430
rect 59782 350 60226 430
rect 60342 350 60786 430
rect 60902 350 61346 430
rect 61462 350 61906 430
rect 62022 350 62466 430
rect 62582 350 63026 430
rect 63142 350 63586 430
rect 63702 350 64146 430
rect 64262 350 64706 430
rect 64822 350 65266 430
rect 65382 350 65826 430
rect 65942 350 66386 430
rect 66502 350 66946 430
rect 67062 350 67506 430
rect 67622 350 68066 430
rect 68182 350 68626 430
rect 68742 350 69186 430
rect 69302 350 69746 430
rect 69862 350 70306 430
rect 70422 350 70866 430
rect 70982 350 71426 430
rect 71542 350 71986 430
rect 72102 350 72546 430
rect 72662 350 73106 430
rect 73222 350 73666 430
rect 73782 350 74226 430
rect 74342 350 74786 430
rect 74902 350 75346 430
rect 75462 350 75906 430
rect 76022 350 76466 430
rect 76582 350 77026 430
rect 77142 350 77586 430
rect 77702 350 78146 430
rect 78262 350 78706 430
rect 78822 350 79266 430
rect 79382 350 79826 430
rect 79942 350 80386 430
rect 80502 350 80946 430
rect 81062 350 81506 430
rect 81622 350 82066 430
rect 82182 350 82626 430
rect 82742 350 83186 430
rect 83302 350 83746 430
rect 83862 350 84306 430
rect 84422 350 84866 430
rect 84982 350 85426 430
rect 85542 350 85986 430
rect 86102 350 86546 430
rect 86662 350 87106 430
rect 87222 350 87666 430
rect 87782 350 88226 430
rect 88342 350 88786 430
rect 88902 350 89346 430
rect 89462 350 89906 430
rect 90022 350 90466 430
rect 90582 350 91026 430
rect 91142 350 91586 430
rect 91702 350 92146 430
rect 92262 350 92706 430
rect 92822 350 93266 430
rect 93382 350 93826 430
rect 93942 350 94386 430
rect 94502 350 94946 430
rect 95062 350 95506 430
rect 95622 350 96066 430
rect 96182 350 96626 430
rect 96742 350 97186 430
rect 97302 350 97746 430
rect 97862 350 98306 430
rect 98422 350 98866 430
rect 98982 350 99426 430
rect 99542 350 99986 430
rect 100102 350 100546 430
rect 100662 350 101106 430
rect 101222 350 101666 430
rect 101782 350 102226 430
rect 102342 350 102786 430
rect 102902 350 103346 430
rect 103462 350 103906 430
rect 104022 350 104466 430
rect 104582 350 105026 430
rect 105142 350 105586 430
rect 105702 350 106146 430
rect 106262 350 106706 430
rect 106822 350 107266 430
rect 107382 350 107826 430
rect 107942 350 108386 430
rect 108502 350 108946 430
rect 109062 350 109506 430
rect 109622 350 110066 430
rect 110182 350 110626 430
rect 110742 350 111186 430
rect 111302 350 111746 430
rect 111862 350 112306 430
rect 112422 350 112866 430
rect 112982 350 113426 430
rect 113542 350 113986 430
rect 114102 350 114546 430
rect 114662 350 115106 430
rect 115222 350 115666 430
rect 115782 350 116226 430
rect 116342 350 116786 430
rect 116902 350 117346 430
rect 117462 350 117906 430
rect 118022 350 118466 430
rect 118582 350 119026 430
rect 119142 350 119586 430
rect 119702 350 120146 430
rect 120262 350 120706 430
rect 120822 350 121266 430
rect 121382 350 121826 430
rect 121942 350 122386 430
rect 122502 350 122946 430
rect 123062 350 123506 430
rect 123622 350 124066 430
rect 124182 350 124626 430
rect 124742 350 125186 430
rect 125302 350 125746 430
rect 125862 350 126306 430
rect 126422 350 126866 430
rect 126982 350 127426 430
rect 127542 350 127986 430
rect 128102 350 128546 430
rect 128662 350 129106 430
rect 129222 350 129666 430
rect 129782 350 130226 430
rect 130342 350 130786 430
rect 130902 350 131346 430
rect 131462 350 131906 430
rect 132022 350 132466 430
rect 132582 350 133026 430
rect 133142 350 133586 430
rect 133702 350 134146 430
rect 134262 350 134706 430
rect 134822 350 135266 430
rect 135382 350 135826 430
rect 135942 350 136386 430
rect 136502 350 136946 430
rect 137062 350 137506 430
rect 137622 350 138066 430
rect 138182 350 138626 430
rect 138742 350 139186 430
rect 139302 350 139746 430
rect 139862 350 140306 430
rect 140422 350 140866 430
rect 140982 350 141426 430
rect 141542 350 141986 430
rect 142102 350 142546 430
rect 142662 350 143106 430
rect 143222 350 143666 430
rect 143782 350 144226 430
rect 144342 350 144786 430
rect 144902 350 145346 430
rect 145462 350 145906 430
rect 146022 350 146466 430
rect 146582 350 147026 430
rect 147142 350 147586 430
rect 147702 350 148146 430
rect 148262 350 148706 430
rect 148822 350 149266 430
rect 149382 350 149826 430
rect 149942 350 150386 430
rect 150502 350 150946 430
rect 151062 350 151506 430
rect 151622 350 152066 430
rect 152182 350 152626 430
rect 152742 350 153186 430
rect 153302 350 153746 430
rect 153862 350 154306 430
rect 154422 350 154866 430
rect 154982 350 155426 430
rect 155542 350 155986 430
rect 156102 350 156546 430
rect 156662 350 157106 430
rect 157222 350 157666 430
rect 157782 350 158226 430
rect 158342 350 158786 430
rect 158902 350 159346 430
rect 159462 350 159906 430
rect 160022 350 160466 430
rect 160582 350 161026 430
rect 161142 350 161586 430
rect 161702 350 162146 430
rect 162262 350 162706 430
rect 162822 350 163266 430
rect 163382 350 163826 430
rect 163942 350 164386 430
rect 164502 350 164946 430
rect 165062 350 165506 430
rect 165622 350 166066 430
rect 166182 350 166626 430
rect 166742 350 167186 430
rect 167302 350 167746 430
rect 167862 350 168306 430
rect 168422 350 168866 430
rect 168982 350 169426 430
rect 169542 350 169986 430
rect 170102 350 170546 430
rect 170662 350 171106 430
rect 171222 350 171666 430
rect 171782 350 172226 430
rect 172342 350 172786 430
rect 172902 350 173346 430
rect 173462 350 173906 430
rect 174022 350 179130 430
<< metal3 >>
rect 0 174944 400 175000
rect 179600 174944 180000 175000
rect 0 167552 400 167608
rect 179600 167552 180000 167608
rect 0 160160 400 160216
rect 179600 160160 180000 160216
rect 0 152768 400 152824
rect 179600 152768 180000 152824
rect 0 145376 400 145432
rect 179600 145376 180000 145432
rect 0 137984 400 138040
rect 179600 137984 180000 138040
rect 0 130592 400 130648
rect 179600 130592 180000 130648
rect 0 123200 400 123256
rect 179600 123200 180000 123256
rect 0 115808 400 115864
rect 179600 115808 180000 115864
rect 0 108416 400 108472
rect 179600 108416 180000 108472
rect 0 101024 400 101080
rect 179600 101024 180000 101080
rect 0 93632 400 93688
rect 179600 93632 180000 93688
rect 0 86240 400 86296
rect 179600 86240 180000 86296
rect 0 78848 400 78904
rect 179600 78848 180000 78904
rect 0 71456 400 71512
rect 179600 71456 180000 71512
rect 0 64064 400 64120
rect 179600 64064 180000 64120
rect 0 56672 400 56728
rect 179600 56672 180000 56728
rect 0 49280 400 49336
rect 179600 49280 180000 49336
rect 0 41888 400 41944
rect 179600 41888 180000 41944
rect 0 34496 400 34552
rect 179600 34496 180000 34552
rect 0 27104 400 27160
rect 179600 27104 180000 27160
rect 0 19712 400 19768
rect 179600 19712 180000 19768
rect 0 12320 400 12376
rect 179600 12320 180000 12376
rect 0 4928 400 4984
rect 179600 4928 180000 4984
<< obsm3 >>
rect 400 175030 179600 178374
rect 430 174914 179570 175030
rect 400 167638 179600 174914
rect 430 167522 179570 167638
rect 400 160246 179600 167522
rect 430 160130 179570 160246
rect 400 152854 179600 160130
rect 430 152738 179570 152854
rect 400 145462 179600 152738
rect 430 145346 179570 145462
rect 400 138070 179600 145346
rect 430 137954 179570 138070
rect 400 130678 179600 137954
rect 430 130562 179570 130678
rect 400 123286 179600 130562
rect 430 123170 179570 123286
rect 400 115894 179600 123170
rect 430 115778 179570 115894
rect 400 108502 179600 115778
rect 430 108386 179570 108502
rect 400 101110 179600 108386
rect 430 100994 179570 101110
rect 400 93718 179600 100994
rect 430 93602 179570 93718
rect 400 86326 179600 93602
rect 430 86210 179570 86326
rect 400 78934 179600 86210
rect 430 78818 179570 78934
rect 400 71542 179600 78818
rect 430 71426 179570 71542
rect 400 64150 179600 71426
rect 430 64034 179570 64150
rect 400 56758 179600 64034
rect 430 56642 179570 56758
rect 400 49366 179600 56642
rect 430 49250 179570 49366
rect 400 41974 179600 49250
rect 430 41858 179570 41974
rect 400 34582 179600 41858
rect 430 34466 179570 34582
rect 400 27190 179600 34466
rect 430 27074 179570 27190
rect 400 19798 179600 27074
rect 430 19682 179570 19798
rect 400 12406 179600 19682
rect 430 12290 179570 12406
rect 400 5014 179600 12290
rect 430 4898 179570 5014
rect 400 518 179600 4898
<< metal4 >>
rect 2224 1538 2384 178390
rect 9904 1538 10064 178390
rect 17584 1538 17744 178390
rect 25264 1538 25424 178390
rect 32944 1538 33104 178390
rect 40624 1538 40784 178390
rect 48304 1538 48464 178390
rect 55984 1538 56144 178390
rect 63664 1538 63824 178390
rect 71344 1538 71504 178390
rect 79024 1538 79184 178390
rect 86704 1538 86864 178390
rect 94384 1538 94544 178390
rect 102064 1538 102224 178390
rect 109744 1538 109904 178390
rect 117424 1538 117584 178390
rect 125104 1538 125264 178390
rect 132784 1538 132944 178390
rect 140464 1538 140624 178390
rect 148144 1538 148304 178390
rect 155824 1538 155984 178390
rect 163504 1538 163664 178390
rect 171184 1538 171344 178390
rect 178864 1538 179024 178390
<< obsm4 >>
rect 3150 1745 9874 175775
rect 10094 1745 17554 175775
rect 17774 1745 25234 175775
rect 25454 1745 32914 175775
rect 33134 1745 40594 175775
rect 40814 1745 48274 175775
rect 48494 1745 55954 175775
rect 56174 1745 63634 175775
rect 63854 1745 71314 175775
rect 71534 1745 78994 175775
rect 79214 1745 86674 175775
rect 86894 1745 94354 175775
rect 94574 1745 102034 175775
rect 102254 1745 109714 175775
rect 109934 1745 117394 175775
rect 117614 1745 125074 175775
rect 125294 1745 132754 175775
rect 132974 1745 140434 175775
rect 140654 1745 148114 175775
rect 148334 1745 155794 175775
rect 156014 1745 163474 175775
rect 163694 1745 171154 175775
rect 171374 1745 174370 175775
<< labels >>
rlabel metal3 s 179600 4928 180000 4984 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 130592 400 130648 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 108416 400 108472 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 86240 400 86296 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 64064 400 64120 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 41888 400 41944 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 19712 400 19768 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 179600 27104 180000 27160 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 179600 49280 180000 49336 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 179600 71456 180000 71512 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 179600 93632 180000 93688 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 179600 115808 180000 115864 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 179600 137984 180000 138040 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 179600 160160 180000 160216 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 174944 400 175000 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 152768 400 152824 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 179600 19712 180000 19768 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 115808 400 115864 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 93632 400 93688 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 71456 400 71512 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 49280 400 49336 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 27104 400 27160 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4928 400 4984 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 179600 41888 180000 41944 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 179600 64064 180000 64120 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 179600 86240 180000 86296 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 179600 108416 180000 108472 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 179600 130592 180000 130648 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 179600 152768 180000 152824 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 179600 174944 180000 175000 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 160160 400 160216 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 137984 400 138040 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 179600 12320 180000 12376 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 123200 400 123256 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 101024 400 101080 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 78848 400 78904 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 56672 400 56728 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 34496 400 34552 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 179600 34496 180000 34552 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 179600 56672 180000 56728 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 179600 78848 180000 78904 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 179600 101024 180000 101080 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 179600 123200 180000 123256 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 179600 145376 180000 145432 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 179600 167552 180000 167608 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 167552 400 167608 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 145376 400 145432 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 172816 0 172872 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 173376 0 173432 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 173936 0 173992 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 65296 0 65352 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 83776 0 83832 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 85456 0 85512 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 87136 0 87192 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 88816 0 88872 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 90496 0 90552 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 92176 0 92232 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 93856 0 93912 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 97216 0 97272 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 98896 0 98952 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 100576 0 100632 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 102256 0 102312 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 103936 0 103992 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 105616 0 105672 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 107296 0 107352 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 110656 0 110712 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 112336 0 112392 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 114016 0 114072 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 117376 0 117432 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 119056 0 119112 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 120736 0 120792 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 122416 0 122472 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 124096 0 124152 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 125776 0 125832 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 127456 0 127512 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 130816 0 130872 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 132496 0 132552 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 134176 0 134232 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 135856 0 135912 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 137536 0 137592 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 139216 0 139272 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 140896 0 140952 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 142576 0 142632 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 144256 0 144312 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 145936 0 145992 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 147616 0 147672 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 72016 0 72072 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 149296 0 149352 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 150976 0 151032 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 152656 0 152712 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 154336 0 154392 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 156016 0 156072 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 157696 0 157752 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 159376 0 159432 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 161056 0 161112 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 162736 0 162792 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 164416 0 164472 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 73696 0 73752 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 166096 0 166152 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 167776 0 167832 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 169456 0 169512 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 171136 0 171192 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 75376 0 75432 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 77056 0 77112 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 78736 0 78792 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 65856 0 65912 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 82656 0 82712 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 84336 0 84392 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 86016 0 86072 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 87696 0 87752 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 89376 0 89432 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 91056 0 91112 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 92736 0 92792 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 94416 0 94472 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 96096 0 96152 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 97776 0 97832 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 99456 0 99512 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 101136 0 101192 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 102816 0 102872 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 104496 0 104552 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 106176 0 106232 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 107856 0 107912 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 109536 0 109592 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 111216 0 111272 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 112896 0 112952 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 114576 0 114632 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 116256 0 116312 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 117936 0 117992 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 119616 0 119672 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 121296 0 121352 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 122976 0 123032 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 124656 0 124712 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 126336 0 126392 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 128016 0 128072 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 129696 0 129752 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 131376 0 131432 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 133056 0 133112 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 134736 0 134792 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 136416 0 136472 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 138096 0 138152 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 139776 0 139832 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 141456 0 141512 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 143136 0 143192 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 144816 0 144872 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 146496 0 146552 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 148176 0 148232 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 72576 0 72632 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 149856 0 149912 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 151536 0 151592 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 153216 0 153272 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 154896 0 154952 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 156576 0 156632 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 158256 0 158312 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 159936 0 159992 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 161616 0 161672 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 163296 0 163352 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 164976 0 165032 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 74256 0 74312 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 166656 0 166712 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 168336 0 168392 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 170016 0 170072 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 171696 0 171752 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 75936 0 75992 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 77616 0 77672 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 79296 0 79352 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 80976 0 81032 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 66416 0 66472 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 83216 0 83272 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 84896 0 84952 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 86576 0 86632 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 88256 0 88312 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 89936 0 89992 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 91616 0 91672 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 94976 0 95032 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 96656 0 96712 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 98336 0 98392 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 100016 0 100072 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 101696 0 101752 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 103376 0 103432 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 105056 0 105112 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 106736 0 106792 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 108416 0 108472 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 110096 0 110152 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 111776 0 111832 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 113456 0 113512 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 115136 0 115192 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 69776 0 69832 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 116816 0 116872 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 118496 0 118552 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 120176 0 120232 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 121856 0 121912 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 123536 0 123592 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 125216 0 125272 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 126896 0 126952 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 128576 0 128632 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 130256 0 130312 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 131936 0 131992 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 133616 0 133672 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 135296 0 135352 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 136976 0 137032 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 138656 0 138712 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 140336 0 140392 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 142016 0 142072 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 143696 0 143752 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 145376 0 145432 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 147056 0 147112 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 148736 0 148792 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 73136 0 73192 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 150416 0 150472 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 152096 0 152152 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 153776 0 153832 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 155456 0 155512 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 157136 0 157192 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 158816 0 158872 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 160496 0 160552 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 162176 0 162232 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 163856 0 163912 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 165536 0 165592 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 74816 0 74872 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 167216 0 167272 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 168896 0 168952 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 170576 0 170632 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 172256 0 172312 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 76496 0 76552 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 78176 0 78232 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 79856 0 79912 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 81536 0 81592 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 178390 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 178390 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 5936 0 5992 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 9296 0 9352 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 36736 0 36792 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 50176 0 50232 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 56896 0 56952 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 58576 0 58632 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 61936 0 61992 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 63616 0 63672 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 40656 0 40712 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 45696 0 45752 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 54096 0 54152 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 55776 0 55832 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 59136 0 59192 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 60816 0 60872 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 29456 0 29512 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 34496 0 34552 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 36176 0 36232 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 41216 0 41272 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 44576 0 44632 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 46256 0 46312 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 47936 0 47992 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 49616 0 49672 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 51296 0 51352 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 52976 0 53032 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 54656 0 54712 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 56336 0 56392 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 59696 0 59752 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 61376 0 61432 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 63056 0 63112 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 64736 0 64792 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 17136 0 17192 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 21056 0 21112 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 22736 0 22792 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 24416 0 24472 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 27776 0 27832 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 10976 0 11032 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 98037494
string GDS_FILE /home/shahid/Desktop/test123/caravel_user_project/openlane/user_proj_example/runs/23_12_07_13_51/results/signoff/user_proj_example.magic.gds
string GDS_START 493242
<< end >>

